`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 19.04.2025 11:06:32
// Design Name: 
// Module Name: mish_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mish_top (
    input  wire [11:0] q57_input,   // 12-bit Q5.7 input
    output wire [31:0] mish_output // 32-bit Q16.16 output
);
    wire [12:0] addr;


    assign addr = q57_input + 13'd2047;

    // Instantiate the ROM module
    mish_rom rom_inst (
        .addr(addr),
        .data_out(mish_output)
    );
endmodule
module mish_rom (
    input  wire [12:0] addr,        // 13-bit address for 8192 entries
    output reg  [31:0] data_out     // 32-bit Q16.16 fixed-point output
);
    // ROM array
    wire [31:0] rom [4095:0];
    assign rom[0]= 32'b00000000000000000000000000000000;
    assign rom[1]= 32'b00000000000000000000000000000000;
    assign rom[2]= 32'b00000000000000000000000000000000;
    assign rom[3]= 32'b00000000000000000000000000000000;
    assign rom[4]= 32'b00000000000000000000000000000000;
    assign rom[5]= 32'b00000000000000000000000000000000;
    assign rom[6]= 32'b00000000000000000000000000000000;
    assign rom[7]= 32'b00000000000000000000000000000000;
    assign rom[8]= 32'b00000000000000000000000000000000;
    assign rom[9]= 32'b00000000000000000000000000000000;
    assign rom[10]= 32'b00000000000000000000000000000000;
    assign rom[11]= 32'b00000000000000000000000000000000;
    assign rom[12]= 32'b00000000000000000000000000000000;
    assign rom[13]= 32'b00000000000000000000000000000000;
    assign rom[14]= 32'b00000000000000000000000000000000;
    assign rom[15]= 32'b00000000000000000000000000000000;
    assign rom[16]= 32'b00000000000000000000000000000000;
    assign rom[17]= 32'b00000000000000000000000000000000;
    assign rom[18]= 32'b00000000000000000000000000000000;
    assign rom[19]= 32'b00000000000000000000000000000000;
    assign rom[20]= 32'b00000000000000000000000000000000;
    assign rom[21]= 32'b00000000000000000000000000000000;
    assign rom[22]= 32'b00000000000000000000000000000000;
    assign rom[23]= 32'b00000000000000000000000000000000;
    assign rom[24]= 32'b00000000000000000000000000000000;
    assign rom[25]= 32'b00000000000000000000000000000000;
    assign rom[26]= 32'b00000000000000000000000000000000;
    assign rom[27]= 32'b00000000000000000000000000000000;
    assign rom[28]= 32'b00000000000000000000000000000000;
    assign rom[29]= 32'b00000000000000000000000000000000;
    assign rom[30]= 32'b00000000000000000000000000000000;
    assign rom[31]= 32'b00000000000000000000000000000000;
    assign rom[32]= 32'b00000000000000000000000000000000;
    assign rom[33]= 32'b00000000000000000000000000000000;
    assign rom[34]= 32'b00000000000000000000000000000000;
    assign rom[35]= 32'b00000000000000000000000000000000;
    assign rom[36]= 32'b00000000000000000000000000000000;
    assign rom[37]= 32'b00000000000000000000000000000000;
    assign rom[38]= 32'b00000000000000000000000000000000;
    assign rom[39]= 32'b00000000000000000000000000000000;
    assign rom[40]= 32'b00000000000000000000000000000000;
    assign rom[41]= 32'b00000000000000000000000000000000;
    assign rom[42]= 32'b00000000000000000000000000000000;
    assign rom[43]= 32'b00000000000000000000000000000000;
    assign rom[44]= 32'b00000000000000000000000000000000;
    assign rom[45]= 32'b00000000000000000000000000000000;
    assign rom[46]= 32'b00000000000000000000000000000000;
    assign rom[47]= 32'b00000000000000000000000000000000;
    assign rom[48]= 32'b00000000000000000000000000000000;
    assign rom[49]= 32'b00000000000000000000000000000000;
    assign rom[50]= 32'b00000000000000000000000000000000;
    assign rom[51]= 32'b00000000000000000000000000000000;
    assign rom[52]= 32'b00000000000000000000000000000000;
    assign rom[53]= 32'b00000000000000000000000000000000;
    assign rom[54]= 32'b00000000000000000000000000000000;
    assign rom[55]= 32'b00000000000000000000000000000000;
    assign rom[56]= 32'b00000000000000000000000000000000;
    assign rom[57]= 32'b00000000000000000000000000000000;
    assign rom[58]= 32'b00000000000000000000000000000000;
    assign rom[59]= 32'b00000000000000000000000000000000;
    assign rom[60]= 32'b00000000000000000000000000000000;
    assign rom[61]= 32'b00000000000000000000000000000000;
    assign rom[62]= 32'b00000000000000000000000000000000;
    assign rom[63]= 32'b00000000000000000000000000000000;
    assign rom[64]= 32'b00000000000000000000000000000000;
    assign rom[65]= 32'b00000000000000000000000000000000;
    assign rom[66]= 32'b00000000000000000000000000000000;
    assign rom[67]= 32'b00000000000000000000000000000000;
    assign rom[68]= 32'b00000000000000000000000000000000;
    assign rom[69]= 32'b00000000000000000000000000000000;
    assign rom[70]= 32'b00000000000000000000000000000000;
    assign rom[71]= 32'b00000000000000000000000000000000;
    assign rom[72]= 32'b00000000000000000000000000000000;
    assign rom[73]= 32'b00000000000000000000000000000000;
    assign rom[74]= 32'b00000000000000000000000000000000;
    assign rom[75]= 32'b00000000000000000000000000000000;
    assign rom[76]= 32'b00000000000000000000000000000000;
    assign rom[77]= 32'b00000000000000000000000000000000;
    assign rom[78]= 32'b00000000000000000000000000000000;
    assign rom[79]= 32'b00000000000000000000000000000000;
    assign rom[80]= 32'b00000000000000000000000000000000;
    assign rom[81]= 32'b00000000000000000000000000000000;
    assign rom[82]= 32'b00000000000000000000000000000000;
    assign rom[83]= 32'b00000000000000000000000000000000;
    assign rom[84]= 32'b00000000000000000000000000000000;
    assign rom[85]= 32'b00000000000000000000000000000000;
    assign rom[86]= 32'b00000000000000000000000000000000;
    assign rom[87]= 32'b00000000000000000000000000000000;
    assign rom[88]= 32'b00000000000000000000000000000000;
    assign rom[89]= 32'b00000000000000000000000000000000;
    assign rom[90]= 32'b00000000000000000000000000000000;
    assign rom[91]= 32'b00000000000000000000000000000000;
    assign rom[92]= 32'b00000000000000000000000000000000;
    assign rom[93]= 32'b00000000000000000000000000000000;
    assign rom[94]= 32'b00000000000000000000000000000000;
    assign rom[95]= 32'b00000000000000000000000000000000;
    assign rom[96]= 32'b00000000000000000000000000000000;
    assign rom[97]= 32'b00000000000000000000000000000000;
    assign rom[98]= 32'b00000000000000000000000000000000;
    assign rom[99]= 32'b00000000000000000000000000000000;
    assign rom[100]= 32'b00000000000000000000000000000000;
    assign rom[101]= 32'b00000000000000000000000000000000;
    assign rom[102]= 32'b00000000000000000000000000000000;
    assign rom[103]= 32'b00000000000000000000000000000000;
    assign rom[104]= 32'b00000000000000000000000000000000;
    assign rom[105]= 32'b00000000000000000000000000000000;
    assign rom[106]= 32'b00000000000000000000000000000000;
    assign rom[107]= 32'b00000000000000000000000000000000;
    assign rom[108]= 32'b00000000000000000000000000000000;
    assign rom[109]= 32'b00000000000000000000000000000000;
    assign rom[110]= 32'b00000000000000000000000000000000;
    assign rom[111]= 32'b00000000000000000000000000000000;
    assign rom[112]= 32'b00000000000000000000000000000000;
    assign rom[113]= 32'b00000000000000000000000000000000;
    assign rom[114]= 32'b00000000000000000000000000000000;
    assign rom[115]= 32'b00000000000000000000000000000000;
    assign rom[116]= 32'b00000000000000000000000000000000;
    assign rom[117]= 32'b00000000000000000000000000000000;
    assign rom[118]= 32'b00000000000000000000000000000000;
    assign rom[119]= 32'b00000000000000000000000000000000;
    assign rom[120]= 32'b00000000000000000000000000000000;
    assign rom[121]= 32'b00000000000000000000000000000000;
    assign rom[122]= 32'b00000000000000000000000000000000;
    assign rom[123]= 32'b00000000000000000000000000000000;
    assign rom[124]= 32'b00000000000000000000000000000000;
    assign rom[125]= 32'b00000000000000000000000000000000;
    assign rom[126]= 32'b00000000000000000000000000000000;
    assign rom[127]= 32'b00000000000000000000000000000000;
    assign rom[128]= 32'b00000000000000000000000000000000;
    assign rom[129]= 32'b00000000000000000000000000000000;
    assign rom[130]= 32'b00000000000000000000000000000000;
    assign rom[131]= 32'b00000000000000000000000000000000;
    assign rom[132]= 32'b00000000000000000000000000000000;
    assign rom[133]= 32'b00000000000000000000000000000000;
    assign rom[134]= 32'b00000000000000000000000000000000;
    assign rom[135]= 32'b00000000000000000000000000000000;
    assign rom[136]= 32'b00000000000000000000000000000000;
    assign rom[137]= 32'b00000000000000000000000000000000;
    assign rom[138]= 32'b00000000000000000000000000000000;
    assign rom[139]= 32'b00000000000000000000000000000000;
    assign rom[140]= 32'b00000000000000000000000000000000;
    assign rom[141]= 32'b00000000000000000000000000000000;
    assign rom[142]= 32'b00000000000000000000000000000000;
    assign rom[143]= 32'b00000000000000000000000000000000;
    assign rom[144]= 32'b00000000000000000000000000000000;
    assign rom[145]= 32'b00000000000000000000000000000000;
    assign rom[146]= 32'b00000000000000000000000000000000;
    assign rom[147]= 32'b00000000000000000000000000000000;
    assign rom[148]= 32'b00000000000000000000000000000000;
    assign rom[149]= 32'b00000000000000000000000000000000;
    assign rom[150]= 32'b00000000000000000000000000000000;
    assign rom[151]= 32'b00000000000000000000000000000000;
    assign rom[152]= 32'b00000000000000000000000000000000;
    assign rom[153]= 32'b00000000000000000000000000000000;
    assign rom[154]= 32'b00000000000000000000000000000000;
    assign rom[155]= 32'b00000000000000000000000000000000;
    assign rom[156]= 32'b00000000000000000000000000000000;
    assign rom[157]= 32'b00000000000000000000000000000000;
    assign rom[158]= 32'b00000000000000000000000000000000;
    assign rom[159]= 32'b00000000000000000000000000000000;
    assign rom[160]= 32'b00000000000000000000000000000000;
    assign rom[161]= 32'b00000000000000000000000000000000;
    assign rom[162]= 32'b00000000000000000000000000000000;
    assign rom[163]= 32'b00000000000000000000000000000000;
    assign rom[164]= 32'b00000000000000000000000000000000;
    assign rom[165]= 32'b00000000000000000000000000000000;
    assign rom[166]= 32'b00000000000000000000000000000000;
    assign rom[167]= 32'b00000000000000000000000000000000;
    assign rom[168]= 32'b00000000000000000000000000000000;
    assign rom[169]= 32'b00000000000000000000000000000000;
    assign rom[170]= 32'b00000000000000000000000000000000;
    assign rom[171]= 32'b00000000000000000000000000000000;
    assign rom[172]= 32'b00000000000000000000000000000000;
    assign rom[173]= 32'b00000000000000000000000000000000;
    assign rom[174]= 32'b00000000000000000000000000000000;
    assign rom[175]= 32'b00000000000000000000000000000000;
    assign rom[176]= 32'b00000000000000000000000000000000;
    assign rom[177]= 32'b00000000000000000000000000000000;
    assign rom[178]= 32'b00000000000000000000000000000000;
    assign rom[179]= 32'b00000000000000000000000000000000;
    assign rom[180]= 32'b00000000000000000000000000000000;
    assign rom[181]= 32'b00000000000000000000000000000000;
    assign rom[182]= 32'b00000000000000000000000000000000;
    assign rom[183]= 32'b00000000000000000000000000000000;
    assign rom[184]= 32'b00000000000000000000000000000000;
    assign rom[185]= 32'b00000000000000000000000000000000;
    assign rom[186]= 32'b00000000000000000000000000000000;
    assign rom[187]= 32'b00000000000000000000000000000000;
    assign rom[188]= 32'b00000000000000000000000000000000;
    assign rom[189]= 32'b00000000000000000000000000000000;
    assign rom[190]= 32'b00000000000000000000000000000000;
    assign rom[191]= 32'b00000000000000000000000000000000;
    assign rom[192]= 32'b00000000000000000000000000000000;
    assign rom[193]= 32'b00000000000000000000000000000000;
    assign rom[194]= 32'b00000000000000000000000000000000;
    assign rom[195]= 32'b00000000000000000000000000000000;
    assign rom[196]= 32'b00000000000000000000000000000000;
    assign rom[197]= 32'b00000000000000000000000000000000;
    assign rom[198]= 32'b00000000000000000000000000000000;
    assign rom[199]= 32'b00000000000000000000000000000000;
    assign rom[200]= 32'b00000000000000000000000000000000;
    assign rom[201]= 32'b00000000000000000000000000000000;
    assign rom[202]= 32'b00000000000000000000000000000000;
    assign rom[203]= 32'b00000000000000000000000000000000;
    assign rom[204]= 32'b00000000000000000000000000000000;
    assign rom[205]= 32'b00000000000000000000000000000000;
    assign rom[206]= 32'b00000000000000000000000000000000;
    assign rom[207]= 32'b00000000000000000000000000000000;
    assign rom[208]= 32'b00000000000000000000000000000000;
    assign rom[209]= 32'b00000000000000000000000000000000;
    assign rom[210]= 32'b00000000000000000000000000000000;
    assign rom[211]= 32'b00000000000000000000000000000000;
    assign rom[212]= 32'b00000000000000000000000000000000;
    assign rom[213]= 32'b00000000000000000000000000000000;
    assign rom[214]= 32'b00000000000000000000000000000000;
    assign rom[215]= 32'b00000000000000000000000000000000;
    assign rom[216]= 32'b00000000000000000000000000000000;
    assign rom[217]= 32'b00000000000000000000000000000000;
    assign rom[218]= 32'b00000000000000000000000000000000;
    assign rom[219]= 32'b00000000000000000000000000000000;
    assign rom[220]= 32'b00000000000000000000000000000000;
    assign rom[221]= 32'b00000000000000000000000000000000;
    assign rom[222]= 32'b00000000000000000000000000000000;
    assign rom[223]= 32'b00000000000000000000000000000000;
    assign rom[224]= 32'b00000000000000000000000000000000;
    assign rom[225]= 32'b00000000000000000000000000000000;
    assign rom[226]= 32'b00000000000000000000000000000000;
    assign rom[227]= 32'b00000000000000000000000000000000;
    assign rom[228]= 32'b00000000000000000000000000000000;
    assign rom[229]= 32'b00000000000000000000000000000000;
    assign rom[230]= 32'b00000000000000000000000000000000;
    assign rom[231]= 32'b00000000000000000000000000000000;
    assign rom[232]= 32'b00000000000000000000000000000000;
    assign rom[233]= 32'b00000000000000000000000000000000;
    assign rom[234]= 32'b00000000000000000000000000000000;
    assign rom[235]= 32'b00000000000000000000000000000000;
    assign rom[236]= 32'b00000000000000000000000000000000;
    assign rom[237]= 32'b00000000000000000000000000000000;
    assign rom[238]= 32'b00000000000000000000000000000000;
    assign rom[239]= 32'b00000000000000000000000000000000;
    assign rom[240]= 32'b00000000000000000000000000000000;
    assign rom[241]= 32'b00000000000000000000000000000000;
    assign rom[242]= 32'b00000000000000000000000000000000;
    assign rom[243]= 32'b00000000000000000000000000000000;
    assign rom[244]= 32'b00000000000000000000000000000000;
    assign rom[245]= 32'b00000000000000000000000000000000;
    assign rom[246]= 32'b00000000000000000000000000000000;
    assign rom[247]= 32'b00000000000000000000000000000000;
    assign rom[248]= 32'b00000000000000000000000000000000;
    assign rom[249]= 32'b00000000000000000000000000000000;
    assign rom[250]= 32'b00000000000000000000000000000000;
    assign rom[251]= 32'b00000000000000000000000000000000;
    assign rom[252]= 32'b00000000000000000000000000000000;
    assign rom[253]= 32'b00000000000000000000000000000000;
    assign rom[254]= 32'b00000000000000000000000000000000;
    assign rom[255]= 32'b00000000000000000000000000000000;
    assign rom[256]= 32'b00000000000000000000000000000000;
    assign rom[257]= 32'b00000000000000000000000000000000;
    assign rom[258]= 32'b00000000000000000000000000000000;
    assign rom[259]= 32'b00000000000000000000000000000000;
    assign rom[260]= 32'b00000000000000000000000000000000;
    assign rom[261]= 32'b00000000000000000000000000000000;
    assign rom[262]= 32'b00000000000000000000000000000000;
    assign rom[263]= 32'b00000000000000000000000000000000;
    assign rom[264]= 32'b00000000000000000000000000000000;
    assign rom[265]= 32'b00000000000000000000000000000000;
    assign rom[266]= 32'b00000000000000000000000000000000;
    assign rom[267]= 32'b00000000000000000000000000000000;
    assign rom[268]= 32'b00000000000000000000000000000000;
    assign rom[269]= 32'b00000000000000000000000000000000;
    assign rom[270]= 32'b00000000000000000000000000000000;
    assign rom[271]= 32'b00000000000000000000000000000000;
    assign rom[272]= 32'b00000000000000000000000000000000;
    assign rom[273]= 32'b00000000000000000000000000000000;
    assign rom[274]= 32'b00000000000000000000000000000000;
    assign rom[275]= 32'b00000000000000000000000000000000;
    assign rom[276]= 32'b00000000000000000000000000000000;
    assign rom[277]= 32'b00000000000000000000000000000000;
    assign rom[278]= 32'b00000000000000000000000000000000;
    assign rom[279]= 32'b00000000000000000000000000000000;
    assign rom[280]= 32'b00000000000000000000000000000000;
    assign rom[281]= 32'b00000000000000000000000000000000;
    assign rom[282]= 32'b00000000000000000000000000000000;
    assign rom[283]= 32'b00000000000000000000000000000000;
    assign rom[284]= 32'b00000000000000000000000000000000;
    assign rom[285]= 32'b00000000000000000000000000000000;
    assign rom[286]= 32'b00000000000000000000000000000000;
    assign rom[287]= 32'b00000000000000000000000000000000;
    assign rom[288]= 32'b00000000000000000000000000000000;
    assign rom[289]= 32'b00000000000000000000000000000000;
    assign rom[290]= 32'b00000000000000000000000000000000;
    assign rom[291]= 32'b00000000000000000000000000000000;
    assign rom[292]= 32'b00000000000000000000000000000000;
    assign rom[293]= 32'b00000000000000000000000000000000;
    assign rom[294]= 32'b11111111111111111111111111111111;
    assign rom[295]= 32'b11111111111111111111111111111111;
    assign rom[296]= 32'b11111111111111111111111111111111;
    assign rom[297]= 32'b11111111111111111111111111111111;
    assign rom[298]= 32'b11111111111111111111111111111111;
    assign rom[299]= 32'b11111111111111111111111111111111;
    assign rom[300]= 32'b11111111111111111111111111111111;
    assign rom[301]= 32'b11111111111111111111111111111111;
    assign rom[302]= 32'b11111111111111111111111111111111;
    assign rom[303]= 32'b11111111111111111111111111111111;
    assign rom[304]= 32'b11111111111111111111111111111111;
    assign rom[305]= 32'b11111111111111111111111111111111;
    assign rom[306]= 32'b11111111111111111111111111111111;
    assign rom[307]= 32'b11111111111111111111111111111111;
    assign rom[308]= 32'b11111111111111111111111111111111;
    assign rom[309]= 32'b11111111111111111111111111111111;
    assign rom[310]= 32'b11111111111111111111111111111111;
    assign rom[311]= 32'b11111111111111111111111111111111;
    assign rom[312]= 32'b11111111111111111111111111111111;
    assign rom[313]= 32'b11111111111111111111111111111111;
    assign rom[314]= 32'b11111111111111111111111111111111;
    assign rom[315]= 32'b11111111111111111111111111111111;
    assign rom[316]= 32'b11111111111111111111111111111111;
    assign rom[317]= 32'b11111111111111111111111111111111;
    assign rom[318]= 32'b11111111111111111111111111111111;
    assign rom[319]= 32'b11111111111111111111111111111111;
    assign rom[320]= 32'b11111111111111111111111111111111;
    assign rom[321]= 32'b11111111111111111111111111111111;
    assign rom[322]= 32'b11111111111111111111111111111111;
    assign rom[323]= 32'b11111111111111111111111111111111;
    assign rom[324]= 32'b11111111111111111111111111111111;
    assign rom[325]= 32'b11111111111111111111111111111111;
    assign rom[326]= 32'b11111111111111111111111111111111;
    assign rom[327]= 32'b11111111111111111111111111111111;
    assign rom[328]= 32'b11111111111111111111111111111111;
    assign rom[329]= 32'b11111111111111111111111111111111;
    assign rom[330]= 32'b11111111111111111111111111111111;
    assign rom[331]= 32'b11111111111111111111111111111111;
    assign rom[332]= 32'b11111111111111111111111111111111;
    assign rom[333]= 32'b11111111111111111111111111111111;
    assign rom[334]= 32'b11111111111111111111111111111111;
    assign rom[335]= 32'b11111111111111111111111111111111;
    assign rom[336]= 32'b11111111111111111111111111111111;
    assign rom[337]= 32'b11111111111111111111111111111111;
    assign rom[338]= 32'b11111111111111111111111111111111;
    assign rom[339]= 32'b11111111111111111111111111111111;
    assign rom[340]= 32'b11111111111111111111111111111111;
    assign rom[341]= 32'b11111111111111111111111111111111;
    assign rom[342]= 32'b11111111111111111111111111111111;
    assign rom[343]= 32'b11111111111111111111111111111111;
    assign rom[344]= 32'b11111111111111111111111111111111;
    assign rom[345]= 32'b11111111111111111111111111111111;
    assign rom[346]= 32'b11111111111111111111111111111111;
    assign rom[347]= 32'b11111111111111111111111111111111;
    assign rom[348]= 32'b11111111111111111111111111111111;
    assign rom[349]= 32'b11111111111111111111111111111111;
    assign rom[350]= 32'b11111111111111111111111111111111;
    assign rom[351]= 32'b11111111111111111111111111111111;
    assign rom[352]= 32'b11111111111111111111111111111111;
    assign rom[353]= 32'b11111111111111111111111111111111;
    assign rom[354]= 32'b11111111111111111111111111111111;
    assign rom[355]= 32'b11111111111111111111111111111111;
    assign rom[356]= 32'b11111111111111111111111111111111;
    assign rom[357]= 32'b11111111111111111111111111111111;
    assign rom[358]= 32'b11111111111111111111111111111111;
    assign rom[359]= 32'b11111111111111111111111111111111;
    assign rom[360]= 32'b11111111111111111111111111111111;
    assign rom[361]= 32'b11111111111111111111111111111111;
    assign rom[362]= 32'b11111111111111111111111111111111;
    assign rom[363]= 32'b11111111111111111111111111111111;
    assign rom[364]= 32'b11111111111111111111111111111111;
    assign rom[365]= 32'b11111111111111111111111111111111;
    assign rom[366]= 32'b11111111111111111111111111111111;
    assign rom[367]= 32'b11111111111111111111111111111111;
    assign rom[368]= 32'b11111111111111111111111111111111;
    assign rom[369]= 32'b11111111111111111111111111111111;
    assign rom[370]= 32'b11111111111111111111111111111111;
    assign rom[371]= 32'b11111111111111111111111111111111;
    assign rom[372]= 32'b11111111111111111111111111111111;
    assign rom[373]= 32'b11111111111111111111111111111111;
    assign rom[374]= 32'b11111111111111111111111111111111;
    assign rom[375]= 32'b11111111111111111111111111111111;
    assign rom[376]= 32'b11111111111111111111111111111111;
    assign rom[377]= 32'b11111111111111111111111111111111;
    assign rom[378]= 32'b11111111111111111111111111111111;
    assign rom[379]= 32'b11111111111111111111111111111111;
    assign rom[380]= 32'b11111111111111111111111111111111;
    assign rom[381]= 32'b11111111111111111111111111111111;
    assign rom[382]= 32'b11111111111111111111111111111111;
    assign rom[383]= 32'b11111111111111111111111111111111;
    assign rom[384]= 32'b11111111111111111111111111111111;
    assign rom[385]= 32'b11111111111111111111111111111111;
    assign rom[386]= 32'b11111111111111111111111111111111;
    assign rom[387]= 32'b11111111111111111111111111111111;
    assign rom[388]= 32'b11111111111111111111111111111111;
    assign rom[389]= 32'b11111111111111111111111111111111;
    assign rom[390]= 32'b11111111111111111111111111111110;
    assign rom[391]= 32'b11111111111111111111111111111110;
    assign rom[392]= 32'b11111111111111111111111111111110;
    assign rom[393]= 32'b11111111111111111111111111111110;
    assign rom[394]= 32'b11111111111111111111111111111110;
    assign rom[395]= 32'b11111111111111111111111111111110;
    assign rom[396]= 32'b11111111111111111111111111111110;
    assign rom[397]= 32'b11111111111111111111111111111110;
    assign rom[398]= 32'b11111111111111111111111111111110;
    assign rom[399]= 32'b11111111111111111111111111111110;
    assign rom[400]= 32'b11111111111111111111111111111110;
    assign rom[401]= 32'b11111111111111111111111111111110;
    assign rom[402]= 32'b11111111111111111111111111111110;
    assign rom[403]= 32'b11111111111111111111111111111110;
    assign rom[404]= 32'b11111111111111111111111111111110;
    assign rom[405]= 32'b11111111111111111111111111111110;
    assign rom[406]= 32'b11111111111111111111111111111110;
    assign rom[407]= 32'b11111111111111111111111111111110;
    assign rom[408]= 32'b11111111111111111111111111111110;
    assign rom[409]= 32'b11111111111111111111111111111110;
    assign rom[410]= 32'b11111111111111111111111111111110;
    assign rom[411]= 32'b11111111111111111111111111111110;
    assign rom[412]= 32'b11111111111111111111111111111110;
    assign rom[413]= 32'b11111111111111111111111111111110;
    assign rom[414]= 32'b11111111111111111111111111111110;
    assign rom[415]= 32'b11111111111111111111111111111110;
    assign rom[416]= 32'b11111111111111111111111111111110;
    assign rom[417]= 32'b11111111111111111111111111111110;
    assign rom[418]= 32'b11111111111111111111111111111110;
    assign rom[419]= 32'b11111111111111111111111111111110;
    assign rom[420]= 32'b11111111111111111111111111111110;
    assign rom[421]= 32'b11111111111111111111111111111110;
    assign rom[422]= 32'b11111111111111111111111111111110;
    assign rom[423]= 32'b11111111111111111111111111111110;
    assign rom[424]= 32'b11111111111111111111111111111110;
    assign rom[425]= 32'b11111111111111111111111111111110;
    assign rom[426]= 32'b11111111111111111111111111111110;
    assign rom[427]= 32'b11111111111111111111111111111110;
    assign rom[428]= 32'b11111111111111111111111111111110;
    assign rom[429]= 32'b11111111111111111111111111111110;
    assign rom[430]= 32'b11111111111111111111111111111110;
    assign rom[431]= 32'b11111111111111111111111111111110;
    assign rom[432]= 32'b11111111111111111111111111111110;
    assign rom[433]= 32'b11111111111111111111111111111110;
    assign rom[434]= 32'b11111111111111111111111111111110;
    assign rom[435]= 32'b11111111111111111111111111111110;
    assign rom[436]= 32'b11111111111111111111111111111110;
    assign rom[437]= 32'b11111111111111111111111111111110;
    assign rom[438]= 32'b11111111111111111111111111111110;
    assign rom[439]= 32'b11111111111111111111111111111110;
    assign rom[440]= 32'b11111111111111111111111111111110;
    assign rom[441]= 32'b11111111111111111111111111111110;
    assign rom[442]= 32'b11111111111111111111111111111110;
    assign rom[443]= 32'b11111111111111111111111111111110;
    assign rom[444]= 32'b11111111111111111111111111111110;
    assign rom[445]= 32'b11111111111111111111111111111110;
    assign rom[446]= 32'b11111111111111111111111111111101;
    assign rom[447]= 32'b11111111111111111111111111111101;
    assign rom[448]= 32'b11111111111111111111111111111101;
    assign rom[449]= 32'b11111111111111111111111111111101;
    assign rom[450]= 32'b11111111111111111111111111111101;
    assign rom[451]= 32'b11111111111111111111111111111101;
    assign rom[452]= 32'b11111111111111111111111111111101;
    assign rom[453]= 32'b11111111111111111111111111111101;
    assign rom[454]= 32'b11111111111111111111111111111101;
    assign rom[455]= 32'b11111111111111111111111111111101;
    assign rom[456]= 32'b11111111111111111111111111111101;
    assign rom[457]= 32'b11111111111111111111111111111101;
    assign rom[458]= 32'b11111111111111111111111111111101;
    assign rom[459]= 32'b11111111111111111111111111111101;
    assign rom[460]= 32'b11111111111111111111111111111101;
    assign rom[461]= 32'b11111111111111111111111111111101;
    assign rom[462]= 32'b11111111111111111111111111111101;
    assign rom[463]= 32'b11111111111111111111111111111101;
    assign rom[464]= 32'b11111111111111111111111111111101;
    assign rom[465]= 32'b11111111111111111111111111111101;
    assign rom[466]= 32'b11111111111111111111111111111101;
    assign rom[467]= 32'b11111111111111111111111111111101;
    assign rom[468]= 32'b11111111111111111111111111111101;
    assign rom[469]= 32'b11111111111111111111111111111101;
    assign rom[470]= 32'b11111111111111111111111111111101;
    assign rom[471]= 32'b11111111111111111111111111111101;
    assign rom[472]= 32'b11111111111111111111111111111101;
    assign rom[473]= 32'b11111111111111111111111111111101;
    assign rom[474]= 32'b11111111111111111111111111111101;
    assign rom[475]= 32'b11111111111111111111111111111101;
    assign rom[476]= 32'b11111111111111111111111111111101;
    assign rom[477]= 32'b11111111111111111111111111111101;
    assign rom[478]= 32'b11111111111111111111111111111101;
    assign rom[479]= 32'b11111111111111111111111111111101;
    assign rom[480]= 32'b11111111111111111111111111111101;
    assign rom[481]= 32'b11111111111111111111111111111101;
    assign rom[482]= 32'b11111111111111111111111111111101;
    assign rom[483]= 32'b11111111111111111111111111111101;
    assign rom[484]= 32'b11111111111111111111111111111101;
    assign rom[485]= 32'b11111111111111111111111111111101;
    assign rom[486]= 32'b11111111111111111111111111111100;
    assign rom[487]= 32'b11111111111111111111111111111100;
    assign rom[488]= 32'b11111111111111111111111111111100;
    assign rom[489]= 32'b11111111111111111111111111111100;
    assign rom[490]= 32'b11111111111111111111111111111100;
    assign rom[491]= 32'b11111111111111111111111111111100;
    assign rom[492]= 32'b11111111111111111111111111111100;
    assign rom[493]= 32'b11111111111111111111111111111100;
    assign rom[494]= 32'b11111111111111111111111111111100;
    assign rom[495]= 32'b11111111111111111111111111111100;
    assign rom[496]= 32'b11111111111111111111111111111100;
    assign rom[497]= 32'b11111111111111111111111111111100;
    assign rom[498]= 32'b11111111111111111111111111111100;
    assign rom[499]= 32'b11111111111111111111111111111100;
    assign rom[500]= 32'b11111111111111111111111111111100;
    assign rom[501]= 32'b11111111111111111111111111111100;
    assign rom[502]= 32'b11111111111111111111111111111100;
    assign rom[503]= 32'b11111111111111111111111111111100;
    assign rom[504]= 32'b11111111111111111111111111111100;
    assign rom[505]= 32'b11111111111111111111111111111100;
    assign rom[506]= 32'b11111111111111111111111111111100;
    assign rom[507]= 32'b11111111111111111111111111111100;
    assign rom[508]= 32'b11111111111111111111111111111100;
    assign rom[509]= 32'b11111111111111111111111111111100;
    assign rom[510]= 32'b11111111111111111111111111111100;
    assign rom[511]= 32'b11111111111111111111111111111100;
    assign rom[512]= 32'b11111111111111111111111111111100;
    assign rom[513]= 32'b11111111111111111111111111111100;
    assign rom[514]= 32'b11111111111111111111111111111100;
    assign rom[515]= 32'b11111111111111111111111111111100;
    assign rom[516]= 32'b11111111111111111111111111111100;
    assign rom[517]= 32'b11111111111111111111111111111011;
    assign rom[518]= 32'b11111111111111111111111111111011;
    assign rom[519]= 32'b11111111111111111111111111111011;
    assign rom[520]= 32'b11111111111111111111111111111011;
    assign rom[521]= 32'b11111111111111111111111111111011;
    assign rom[522]= 32'b11111111111111111111111111111011;
    assign rom[523]= 32'b11111111111111111111111111111011;
    assign rom[524]= 32'b11111111111111111111111111111011;
    assign rom[525]= 32'b11111111111111111111111111111011;
    assign rom[526]= 32'b11111111111111111111111111111011;
    assign rom[527]= 32'b11111111111111111111111111111011;
    assign rom[528]= 32'b11111111111111111111111111111011;
    assign rom[529]= 32'b11111111111111111111111111111011;
    assign rom[530]= 32'b11111111111111111111111111111011;
    assign rom[531]= 32'b11111111111111111111111111111011;
    assign rom[532]= 32'b11111111111111111111111111111011;
    assign rom[533]= 32'b11111111111111111111111111111011;
    assign rom[534]= 32'b11111111111111111111111111111011;
    assign rom[535]= 32'b11111111111111111111111111111011;
    assign rom[536]= 32'b11111111111111111111111111111011;
    assign rom[537]= 32'b11111111111111111111111111111011;
    assign rom[538]= 32'b11111111111111111111111111111011;
    assign rom[539]= 32'b11111111111111111111111111111011;
    assign rom[540]= 32'b11111111111111111111111111111011;
    assign rom[541]= 32'b11111111111111111111111111111011;
    assign rom[542]= 32'b11111111111111111111111111111011;
    assign rom[543]= 32'b11111111111111111111111111111010;
    assign rom[544]= 32'b11111111111111111111111111111010;
    assign rom[545]= 32'b11111111111111111111111111111010;
    assign rom[546]= 32'b11111111111111111111111111111010;
    assign rom[547]= 32'b11111111111111111111111111111010;
    assign rom[548]= 32'b11111111111111111111111111111010;
    assign rom[549]= 32'b11111111111111111111111111111010;
    assign rom[550]= 32'b11111111111111111111111111111010;
    assign rom[551]= 32'b11111111111111111111111111111010;
    assign rom[552]= 32'b11111111111111111111111111111010;
    assign rom[553]= 32'b11111111111111111111111111111010;
    assign rom[554]= 32'b11111111111111111111111111111010;
    assign rom[555]= 32'b11111111111111111111111111111010;
    assign rom[556]= 32'b11111111111111111111111111111010;
    assign rom[557]= 32'b11111111111111111111111111111010;
    assign rom[558]= 32'b11111111111111111111111111111010;
    assign rom[559]= 32'b11111111111111111111111111111010;
    assign rom[560]= 32'b11111111111111111111111111111010;
    assign rom[561]= 32'b11111111111111111111111111111010;
    assign rom[562]= 32'b11111111111111111111111111111010;
    assign rom[563]= 32'b11111111111111111111111111111010;
    assign rom[564]= 32'b11111111111111111111111111111001;
    assign rom[565]= 32'b11111111111111111111111111111001;
    assign rom[566]= 32'b11111111111111111111111111111001;
    assign rom[567]= 32'b11111111111111111111111111111001;
    assign rom[568]= 32'b11111111111111111111111111111001;
    assign rom[569]= 32'b11111111111111111111111111111001;
    assign rom[570]= 32'b11111111111111111111111111111001;
    assign rom[571]= 32'b11111111111111111111111111111001;
    assign rom[572]= 32'b11111111111111111111111111111001;
    assign rom[573]= 32'b11111111111111111111111111111001;
    assign rom[574]= 32'b11111111111111111111111111111001;
    assign rom[575]= 32'b11111111111111111111111111111001;
    assign rom[576]= 32'b11111111111111111111111111111001;
    assign rom[577]= 32'b11111111111111111111111111111001;
    assign rom[578]= 32'b11111111111111111111111111111001;
    assign rom[579]= 32'b11111111111111111111111111111001;
    assign rom[580]= 32'b11111111111111111111111111111001;
    assign rom[581]= 32'b11111111111111111111111111111001;
    assign rom[582]= 32'b11111111111111111111111111111001;
    assign rom[583]= 32'b11111111111111111111111111111000;
    assign rom[584]= 32'b11111111111111111111111111111000;
    assign rom[585]= 32'b11111111111111111111111111111000;
    assign rom[586]= 32'b11111111111111111111111111111000;
    assign rom[587]= 32'b11111111111111111111111111111000;
    assign rom[588]= 32'b11111111111111111111111111111000;
    assign rom[589]= 32'b11111111111111111111111111111000;
    assign rom[590]= 32'b11111111111111111111111111111000;
    assign rom[591]= 32'b11111111111111111111111111111000;
    assign rom[592]= 32'b11111111111111111111111111111000;
    assign rom[593]= 32'b11111111111111111111111111111000;
    assign rom[594]= 32'b11111111111111111111111111111000;
    assign rom[595]= 32'b11111111111111111111111111111000;
    assign rom[596]= 32'b11111111111111111111111111111000;
    assign rom[597]= 32'b11111111111111111111111111111000;
    assign rom[598]= 32'b11111111111111111111111111111000;
    assign rom[599]= 32'b11111111111111111111111111111000;
    assign rom[600]= 32'b11111111111111111111111111110111;
    assign rom[601]= 32'b11111111111111111111111111110111;
    assign rom[602]= 32'b11111111111111111111111111110111;
    assign rom[603]= 32'b11111111111111111111111111110111;
    assign rom[604]= 32'b11111111111111111111111111110111;
    assign rom[605]= 32'b11111111111111111111111111110111;
    assign rom[606]= 32'b11111111111111111111111111110111;
    assign rom[607]= 32'b11111111111111111111111111110111;
    assign rom[608]= 32'b11111111111111111111111111110111;
    assign rom[609]= 32'b11111111111111111111111111110111;
    assign rom[610]= 32'b11111111111111111111111111110111;
    assign rom[611]= 32'b11111111111111111111111111110111;
    assign rom[612]= 32'b11111111111111111111111111110111;
    assign rom[613]= 32'b11111111111111111111111111110111;
    assign rom[614]= 32'b11111111111111111111111111110110;
    assign rom[615]= 32'b11111111111111111111111111110110;
    assign rom[616]= 32'b11111111111111111111111111110110;
    assign rom[617]= 32'b11111111111111111111111111110110;
    assign rom[618]= 32'b11111111111111111111111111110110;
    assign rom[619]= 32'b11111111111111111111111111110110;
    assign rom[620]= 32'b11111111111111111111111111110110;
    assign rom[621]= 32'b11111111111111111111111111110110;
    assign rom[622]= 32'b11111111111111111111111111110110;
    assign rom[623]= 32'b11111111111111111111111111110110;
    assign rom[624]= 32'b11111111111111111111111111110110;
    assign rom[625]= 32'b11111111111111111111111111110110;
    assign rom[626]= 32'b11111111111111111111111111110110;
    assign rom[627]= 32'b11111111111111111111111111110110;
    assign rom[628]= 32'b11111111111111111111111111110101;
    assign rom[629]= 32'b11111111111111111111111111110101;
    assign rom[630]= 32'b11111111111111111111111111110101;
    assign rom[631]= 32'b11111111111111111111111111110101;
    assign rom[632]= 32'b11111111111111111111111111110101;
    assign rom[633]= 32'b11111111111111111111111111110101;
    assign rom[634]= 32'b11111111111111111111111111110101;
    assign rom[635]= 32'b11111111111111111111111111110101;
    assign rom[636]= 32'b11111111111111111111111111110101;
    assign rom[637]= 32'b11111111111111111111111111110101;
    assign rom[638]= 32'b11111111111111111111111111110101;
    assign rom[639]= 32'b11111111111111111111111111110101;
    assign rom[640]= 32'b11111111111111111111111111110100;
    assign rom[641]= 32'b11111111111111111111111111110100;
    assign rom[642]= 32'b11111111111111111111111111110100;
    assign rom[643]= 32'b11111111111111111111111111110100;
    assign rom[644]= 32'b11111111111111111111111111110100;
    assign rom[645]= 32'b11111111111111111111111111110100;
    assign rom[646]= 32'b11111111111111111111111111110100;
    assign rom[647]= 32'b11111111111111111111111111110100;
    assign rom[648]= 32'b11111111111111111111111111110100;
    assign rom[649]= 32'b11111111111111111111111111110100;
    assign rom[650]= 32'b11111111111111111111111111110100;
    assign rom[651]= 32'b11111111111111111111111111110011;
    assign rom[652]= 32'b11111111111111111111111111110011;
    assign rom[653]= 32'b11111111111111111111111111110011;
    assign rom[654]= 32'b11111111111111111111111111110011;
    assign rom[655]= 32'b11111111111111111111111111110011;
    assign rom[656]= 32'b11111111111111111111111111110011;
    assign rom[657]= 32'b11111111111111111111111111110011;
    assign rom[658]= 32'b11111111111111111111111111110011;
    assign rom[659]= 32'b11111111111111111111111111110011;
    assign rom[660]= 32'b11111111111111111111111111110011;
    assign rom[661]= 32'b11111111111111111111111111110011;
    assign rom[662]= 32'b11111111111111111111111111110010;
    assign rom[663]= 32'b11111111111111111111111111110010;
    assign rom[664]= 32'b11111111111111111111111111110010;
    assign rom[665]= 32'b11111111111111111111111111110010;
    assign rom[666]= 32'b11111111111111111111111111110010;
    assign rom[667]= 32'b11111111111111111111111111110010;
    assign rom[668]= 32'b11111111111111111111111111110010;
    assign rom[669]= 32'b11111111111111111111111111110010;
    assign rom[670]= 32'b11111111111111111111111111110010;
    assign rom[671]= 32'b11111111111111111111111111110001;
    assign rom[672]= 32'b11111111111111111111111111110001;
    assign rom[673]= 32'b11111111111111111111111111110001;
    assign rom[674]= 32'b11111111111111111111111111110001;
    assign rom[675]= 32'b11111111111111111111111111110001;
    assign rom[676]= 32'b11111111111111111111111111110001;
    assign rom[677]= 32'b11111111111111111111111111110001;
    assign rom[678]= 32'b11111111111111111111111111110001;
    assign rom[679]= 32'b11111111111111111111111111110001;
    assign rom[680]= 32'b11111111111111111111111111110001;
    assign rom[681]= 32'b11111111111111111111111111110000;
    assign rom[682]= 32'b11111111111111111111111111110000;
    assign rom[683]= 32'b11111111111111111111111111110000;
    assign rom[684]= 32'b11111111111111111111111111110000;
    assign rom[685]= 32'b11111111111111111111111111110000;
    assign rom[686]= 32'b11111111111111111111111111110000;
    assign rom[687]= 32'b11111111111111111111111111110000;
    assign rom[688]= 32'b11111111111111111111111111110000;
    assign rom[689]= 32'b11111111111111111111111111101111;
    assign rom[690]= 32'b11111111111111111111111111101111;
    assign rom[691]= 32'b11111111111111111111111111101111;
    assign rom[692]= 32'b11111111111111111111111111101111;
    assign rom[693]= 32'b11111111111111111111111111101111;
    assign rom[694]= 32'b11111111111111111111111111101111;
    assign rom[695]= 32'b11111111111111111111111111101111;
    assign rom[696]= 32'b11111111111111111111111111101111;
    assign rom[697]= 32'b11111111111111111111111111101110;
    assign rom[698]= 32'b11111111111111111111111111101110;
    assign rom[699]= 32'b11111111111111111111111111101110;
    assign rom[700]= 32'b11111111111111111111111111101110;
    assign rom[701]= 32'b11111111111111111111111111101110;
    assign rom[702]= 32'b11111111111111111111111111101110;
    assign rom[703]= 32'b11111111111111111111111111101110;
    assign rom[704]= 32'b11111111111111111111111111101110;
    assign rom[705]= 32'b11111111111111111111111111101101;
    assign rom[706]= 32'b11111111111111111111111111101101;
    assign rom[707]= 32'b11111111111111111111111111101101;
    assign rom[708]= 32'b11111111111111111111111111101101;
    assign rom[709]= 32'b11111111111111111111111111101101;
    assign rom[710]= 32'b11111111111111111111111111101101;
    assign rom[711]= 32'b11111111111111111111111111101101;
    assign rom[712]= 32'b11111111111111111111111111101100;
    assign rom[713]= 32'b11111111111111111111111111101100;
    assign rom[714]= 32'b11111111111111111111111111101100;
    assign rom[715]= 32'b11111111111111111111111111101100;
    assign rom[716]= 32'b11111111111111111111111111101100;
    assign rom[717]= 32'b11111111111111111111111111101100;
    assign rom[718]= 32'b11111111111111111111111111101100;
    assign rom[719]= 32'b11111111111111111111111111101011;
    assign rom[720]= 32'b11111111111111111111111111101011;
    assign rom[721]= 32'b11111111111111111111111111101011;
    assign rom[722]= 32'b11111111111111111111111111101011;
    assign rom[723]= 32'b11111111111111111111111111101011;
    assign rom[724]= 32'b11111111111111111111111111101011;
    assign rom[725]= 32'b11111111111111111111111111101011;
    assign rom[726]= 32'b11111111111111111111111111101010;
    assign rom[727]= 32'b11111111111111111111111111101010;
    assign rom[728]= 32'b11111111111111111111111111101010;
    assign rom[729]= 32'b11111111111111111111111111101010;
    assign rom[730]= 32'b11111111111111111111111111101010;
    assign rom[731]= 32'b11111111111111111111111111101010;
    assign rom[732]= 32'b11111111111111111111111111101001;
    assign rom[733]= 32'b11111111111111111111111111101001;
    assign rom[734]= 32'b11111111111111111111111111101001;
    assign rom[735]= 32'b11111111111111111111111111101001;
    assign rom[736]= 32'b11111111111111111111111111101001;
    assign rom[737]= 32'b11111111111111111111111111101001;
    assign rom[738]= 32'b11111111111111111111111111101000;
    assign rom[739]= 32'b11111111111111111111111111101000;
    assign rom[740]= 32'b11111111111111111111111111101000;
    assign rom[741]= 32'b11111111111111111111111111101000;
    assign rom[742]= 32'b11111111111111111111111111101000;
    assign rom[743]= 32'b11111111111111111111111111101000;
    assign rom[744]= 32'b11111111111111111111111111100111;
    assign rom[745]= 32'b11111111111111111111111111100111;
    assign rom[746]= 32'b11111111111111111111111111100111;
    assign rom[747]= 32'b11111111111111111111111111100111;
    assign rom[748]= 32'b11111111111111111111111111100111;
    assign rom[749]= 32'b11111111111111111111111111100110;
    assign rom[750]= 32'b11111111111111111111111111100110;
    assign rom[751]= 32'b11111111111111111111111111100110;
    assign rom[752]= 32'b11111111111111111111111111100110;
    assign rom[753]= 32'b11111111111111111111111111100110;
    assign rom[754]= 32'b11111111111111111111111111100110;
    assign rom[755]= 32'b11111111111111111111111111100101;
    assign rom[756]= 32'b11111111111111111111111111100101;
    assign rom[757]= 32'b11111111111111111111111111100101;
    assign rom[758]= 32'b11111111111111111111111111100101;
    assign rom[759]= 32'b11111111111111111111111111100101;
    assign rom[760]= 32'b11111111111111111111111111100100;
    assign rom[761]= 32'b11111111111111111111111111100100;
    assign rom[762]= 32'b11111111111111111111111111100100;
    assign rom[763]= 32'b11111111111111111111111111100100;
    assign rom[764]= 32'b11111111111111111111111111100100;
    assign rom[765]= 32'b11111111111111111111111111100011;
    assign rom[766]= 32'b11111111111111111111111111100011;
    assign rom[767]= 32'b11111111111111111111111111100011;
    assign rom[768]= 32'b11111111111111111111111111100011;
    assign rom[769]= 32'b11111111111111111111111111100011;
    assign rom[770]= 32'b11111111111111111111111111100010;
    assign rom[771]= 32'b11111111111111111111111111100010;
    assign rom[772]= 32'b11111111111111111111111111100010;
    assign rom[773]= 32'b11111111111111111111111111100010;
    assign rom[774]= 32'b11111111111111111111111111100001;
    assign rom[775]= 32'b11111111111111111111111111100001;
    assign rom[776]= 32'b11111111111111111111111111100001;
    assign rom[777]= 32'b11111111111111111111111111100001;
    assign rom[778]= 32'b11111111111111111111111111100001;
    assign rom[779]= 32'b11111111111111111111111111100000;
    assign rom[780]= 32'b11111111111111111111111111100000;
    assign rom[781]= 32'b11111111111111111111111111100000;
    assign rom[782]= 32'b11111111111111111111111111100000;
    assign rom[783]= 32'b11111111111111111111111111011111;
    assign rom[784]= 32'b11111111111111111111111111011111;
    assign rom[785]= 32'b11111111111111111111111111011111;
    assign rom[786]= 32'b11111111111111111111111111011111;
    assign rom[787]= 32'b11111111111111111111111111011110;
    assign rom[788]= 32'b11111111111111111111111111011110;
    assign rom[789]= 32'b11111111111111111111111111011110;
    assign rom[790]= 32'b11111111111111111111111111011110;
    assign rom[791]= 32'b11111111111111111111111111011110;
    assign rom[792]= 32'b11111111111111111111111111011101;
    assign rom[793]= 32'b11111111111111111111111111011101;
    assign rom[794]= 32'b11111111111111111111111111011101;
    assign rom[795]= 32'b11111111111111111111111111011101;
    assign rom[796]= 32'b11111111111111111111111111011100;
    assign rom[797]= 32'b11111111111111111111111111011100;
    assign rom[798]= 32'b11111111111111111111111111011100;
    assign rom[799]= 32'b11111111111111111111111111011100;
    assign rom[800]= 32'b11111111111111111111111111011011;
    assign rom[801]= 32'b11111111111111111111111111011011;
    assign rom[802]= 32'b11111111111111111111111111011011;
    assign rom[803]= 32'b11111111111111111111111111011010;
    assign rom[804]= 32'b11111111111111111111111111011010;
    assign rom[805]= 32'b11111111111111111111111111011010;
    assign rom[806]= 32'b11111111111111111111111111011010;
    assign rom[807]= 32'b11111111111111111111111111011001;
    assign rom[808]= 32'b11111111111111111111111111011001;
    assign rom[809]= 32'b11111111111111111111111111011001;
    assign rom[810]= 32'b11111111111111111111111111011001;
    assign rom[811]= 32'b11111111111111111111111111011000;
    assign rom[812]= 32'b11111111111111111111111111011000;
    assign rom[813]= 32'b11111111111111111111111111011000;
    assign rom[814]= 32'b11111111111111111111111111010111;
    assign rom[815]= 32'b11111111111111111111111111010111;
    assign rom[816]= 32'b11111111111111111111111111010111;
    assign rom[817]= 32'b11111111111111111111111111010111;
    assign rom[818]= 32'b11111111111111111111111111010110;
    assign rom[819]= 32'b11111111111111111111111111010110;
    assign rom[820]= 32'b11111111111111111111111111010110;
    assign rom[821]= 32'b11111111111111111111111111010101;
    assign rom[822]= 32'b11111111111111111111111111010101;
    assign rom[823]= 32'b11111111111111111111111111010101;
    assign rom[824]= 32'b11111111111111111111111111010100;
    assign rom[825]= 32'b11111111111111111111111111010100;
    assign rom[826]= 32'b11111111111111111111111111010100;
    assign rom[827]= 32'b11111111111111111111111111010100;
    assign rom[828]= 32'b11111111111111111111111111010011;
    assign rom[829]= 32'b11111111111111111111111111010011;
    assign rom[830]= 32'b11111111111111111111111111010011;
    assign rom[831]= 32'b11111111111111111111111111010010;
    assign rom[832]= 32'b11111111111111111111111111010010;
    assign rom[833]= 32'b11111111111111111111111111010010;
    assign rom[834]= 32'b11111111111111111111111111010001;
    assign rom[835]= 32'b11111111111111111111111111010001;
    assign rom[836]= 32'b11111111111111111111111111010001;
    assign rom[837]= 32'b11111111111111111111111111010000;
    assign rom[838]= 32'b11111111111111111111111111010000;
    assign rom[839]= 32'b11111111111111111111111111010000;
    assign rom[840]= 32'b11111111111111111111111111001111;
    assign rom[841]= 32'b11111111111111111111111111001111;
    assign rom[842]= 32'b11111111111111111111111111001111;
    assign rom[843]= 32'b11111111111111111111111111001110;
    assign rom[844]= 32'b11111111111111111111111111001110;
    assign rom[845]= 32'b11111111111111111111111111001101;
    assign rom[846]= 32'b11111111111111111111111111001101;
    assign rom[847]= 32'b11111111111111111111111111001101;
    assign rom[848]= 32'b11111111111111111111111111001100;
    assign rom[849]= 32'b11111111111111111111111111001100;
    assign rom[850]= 32'b11111111111111111111111111001100;
    assign rom[851]= 32'b11111111111111111111111111001011;
    assign rom[852]= 32'b11111111111111111111111111001011;
    assign rom[853]= 32'b11111111111111111111111111001011;
    assign rom[854]= 32'b11111111111111111111111111001010;
    assign rom[855]= 32'b11111111111111111111111111001010;
    assign rom[856]= 32'b11111111111111111111111111001001;
    assign rom[857]= 32'b11111111111111111111111111001001;
    assign rom[858]= 32'b11111111111111111111111111001001;
    assign rom[859]= 32'b11111111111111111111111111001000;
    assign rom[860]= 32'b11111111111111111111111111001000;
    assign rom[861]= 32'b11111111111111111111111111000111;
    assign rom[862]= 32'b11111111111111111111111111000111;
    assign rom[863]= 32'b11111111111111111111111111000111;
    assign rom[864]= 32'b11111111111111111111111111000110;
    assign rom[865]= 32'b11111111111111111111111111000110;
    assign rom[866]= 32'b11111111111111111111111111000101;
    assign rom[867]= 32'b11111111111111111111111111000101;
    assign rom[868]= 32'b11111111111111111111111111000101;
    assign rom[869]= 32'b11111111111111111111111111000100;
    assign rom[870]= 32'b11111111111111111111111111000100;
    assign rom[871]= 32'b11111111111111111111111111000011;
    assign rom[872]= 32'b11111111111111111111111111000011;
    assign rom[873]= 32'b11111111111111111111111111000010;
    assign rom[874]= 32'b11111111111111111111111111000010;
    assign rom[875]= 32'b11111111111111111111111111000010;
    assign rom[876]= 32'b11111111111111111111111111000001;
    assign rom[877]= 32'b11111111111111111111111111000001;
    assign rom[878]= 32'b11111111111111111111111111000000;
    assign rom[879]= 32'b11111111111111111111111111000000;
    assign rom[880]= 32'b11111111111111111111111110111111;
    assign rom[881]= 32'b11111111111111111111111110111111;
    assign rom[882]= 32'b11111111111111111111111110111110;
    assign rom[883]= 32'b11111111111111111111111110111110;
    assign rom[884]= 32'b11111111111111111111111110111110;
    assign rom[885]= 32'b11111111111111111111111110111101;
    assign rom[886]= 32'b11111111111111111111111110111101;
    assign rom[887]= 32'b11111111111111111111111110111100;
    assign rom[888]= 32'b11111111111111111111111110111100;
    assign rom[889]= 32'b11111111111111111111111110111011;
    assign rom[890]= 32'b11111111111111111111111110111011;
    assign rom[891]= 32'b11111111111111111111111110111010;
    assign rom[892]= 32'b11111111111111111111111110111010;
    assign rom[893]= 32'b11111111111111111111111110111001;
    assign rom[894]= 32'b11111111111111111111111110111001;
    assign rom[895]= 32'b11111111111111111111111110111000;
    assign rom[896]= 32'b11111111111111111111111110111000;
    assign rom[897]= 32'b11111111111111111111111110110111;
    assign rom[898]= 32'b11111111111111111111111110110111;
    assign rom[899]= 32'b11111111111111111111111110110110;
    assign rom[900]= 32'b11111111111111111111111110110110;
    assign rom[901]= 32'b11111111111111111111111110110101;
    assign rom[902]= 32'b11111111111111111111111110110101;
    assign rom[903]= 32'b11111111111111111111111110110100;
    assign rom[904]= 32'b11111111111111111111111110110100;
    assign rom[905]= 32'b11111111111111111111111110110011;
    assign rom[906]= 32'b11111111111111111111111110110010;
    assign rom[907]= 32'b11111111111111111111111110110010;
    assign rom[908]= 32'b11111111111111111111111110110001;
    assign rom[909]= 32'b11111111111111111111111110110001;
    assign rom[910]= 32'b11111111111111111111111110110000;
    assign rom[911]= 32'b11111111111111111111111110110000;
    assign rom[912]= 32'b11111111111111111111111110101111;
    assign rom[913]= 32'b11111111111111111111111110101111;
    assign rom[914]= 32'b11111111111111111111111110101110;
    assign rom[915]= 32'b11111111111111111111111110101101;
    assign rom[916]= 32'b11111111111111111111111110101101;
    assign rom[917]= 32'b11111111111111111111111110101100;
    assign rom[918]= 32'b11111111111111111111111110101100;
    assign rom[919]= 32'b11111111111111111111111110101011;
    assign rom[920]= 32'b11111111111111111111111110101011;
    assign rom[921]= 32'b11111111111111111111111110101010;
    assign rom[922]= 32'b11111111111111111111111110101001;
    assign rom[923]= 32'b11111111111111111111111110101001;
    assign rom[924]= 32'b11111111111111111111111110101000;
    assign rom[925]= 32'b11111111111111111111111110101000;
    assign rom[926]= 32'b11111111111111111111111110100111;
    assign rom[927]= 32'b11111111111111111111111110100110;
    assign rom[928]= 32'b11111111111111111111111110100110;
    assign rom[929]= 32'b11111111111111111111111110100101;
    assign rom[930]= 32'b11111111111111111111111110100100;
    assign rom[931]= 32'b11111111111111111111111110100100;
    assign rom[932]= 32'b11111111111111111111111110100011;
    assign rom[933]= 32'b11111111111111111111111110100010;
    assign rom[934]= 32'b11111111111111111111111110100010;
    assign rom[935]= 32'b11111111111111111111111110100001;
    assign rom[936]= 32'b11111111111111111111111110100000;
    assign rom[937]= 32'b11111111111111111111111110100000;
    assign rom[938]= 32'b11111111111111111111111110011111;
    assign rom[939]= 32'b11111111111111111111111110011110;
    assign rom[940]= 32'b11111111111111111111111110011110;
    assign rom[941]= 32'b11111111111111111111111110011101;
    assign rom[942]= 32'b11111111111111111111111110011100;
    assign rom[943]= 32'b11111111111111111111111110011100;
    assign rom[944]= 32'b11111111111111111111111110011011;
    assign rom[945]= 32'b11111111111111111111111110011010;
    assign rom[946]= 32'b11111111111111111111111110011010;
    assign rom[947]= 32'b11111111111111111111111110011001;
    assign rom[948]= 32'b11111111111111111111111110011000;
    assign rom[949]= 32'b11111111111111111111111110010111;
    assign rom[950]= 32'b11111111111111111111111110010111;
    assign rom[951]= 32'b11111111111111111111111110010110;
    assign rom[952]= 32'b11111111111111111111111110010101;
    assign rom[953]= 32'b11111111111111111111111110010101;
    assign rom[954]= 32'b11111111111111111111111110010100;
    assign rom[955]= 32'b11111111111111111111111110010011;
    assign rom[956]= 32'b11111111111111111111111110010010;
    assign rom[957]= 32'b11111111111111111111111110010001;
    assign rom[958]= 32'b11111111111111111111111110010001;
    assign rom[959]= 32'b11111111111111111111111110010000;
    assign rom[960]= 32'b11111111111111111111111110001111;
    assign rom[961]= 32'b11111111111111111111111110001110;
    assign rom[962]= 32'b11111111111111111111111110001110;
    assign rom[963]= 32'b11111111111111111111111110001101;
    assign rom[964]= 32'b11111111111111111111111110001100;
    assign rom[965]= 32'b11111111111111111111111110001011;
    assign rom[966]= 32'b11111111111111111111111110001010;
    assign rom[967]= 32'b11111111111111111111111110001010;
    assign rom[968]= 32'b11111111111111111111111110001001;
    assign rom[969]= 32'b11111111111111111111111110001000;
    assign rom[970]= 32'b11111111111111111111111110000111;
    assign rom[971]= 32'b11111111111111111111111110000110;
    assign rom[972]= 32'b11111111111111111111111110000101;
    assign rom[973]= 32'b11111111111111111111111110000101;
    assign rom[974]= 32'b11111111111111111111111110000100;
    assign rom[975]= 32'b11111111111111111111111110000011;
    assign rom[976]= 32'b11111111111111111111111110000010;
    assign rom[977]= 32'b11111111111111111111111110000001;
    assign rom[978]= 32'b11111111111111111111111110000000;
    assign rom[979]= 32'b11111111111111111111111101111111;
    assign rom[980]= 32'b11111111111111111111111101111110;
    assign rom[981]= 32'b11111111111111111111111101111110;
    assign rom[982]= 32'b11111111111111111111111101111101;
    assign rom[983]= 32'b11111111111111111111111101111100;
    assign rom[984]= 32'b11111111111111111111111101111011;
    assign rom[985]= 32'b11111111111111111111111101111010;
    assign rom[986]= 32'b11111111111111111111111101111001;
    assign rom[987]= 32'b11111111111111111111111101111000;
    assign rom[988]= 32'b11111111111111111111111101110111;
    assign rom[989]= 32'b11111111111111111111111101110110;
    assign rom[990]= 32'b11111111111111111111111101110101;
    assign rom[991]= 32'b11111111111111111111111101110100;
    assign rom[992]= 32'b11111111111111111111111101110011;
    assign rom[993]= 32'b11111111111111111111111101110010;
    assign rom[994]= 32'b11111111111111111111111101110001;
    assign rom[995]= 32'b11111111111111111111111101110000;
    assign rom[996]= 32'b11111111111111111111111101101111;
    assign rom[997]= 32'b11111111111111111111111101101110;
    assign rom[998]= 32'b11111111111111111111111101101101;
    assign rom[999]= 32'b11111111111111111111111101101100;
    assign rom[1000]= 32'b11111111111111111111111101101011;
    assign rom[1001]= 32'b11111111111111111111111101101010;
    assign rom[1002]= 32'b11111111111111111111111101101001;
    assign rom[1003]= 32'b11111111111111111111111101101000;
    assign rom[1004]= 32'b11111111111111111111111101100111;
    assign rom[1005]= 32'b11111111111111111111111101100110;
    assign rom[1006]= 32'b11111111111111111111111101100101;
    assign rom[1007]= 32'b11111111111111111111111101100100;
    assign rom[1008]= 32'b11111111111111111111111101100011;
    assign rom[1009]= 32'b11111111111111111111111101100010;
    assign rom[1010]= 32'b11111111111111111111111101100001;
    assign rom[1011]= 32'b11111111111111111111111101100000;
    assign rom[1012]= 32'b11111111111111111111111101011111;
    assign rom[1013]= 32'b11111111111111111111111101011101;
    assign rom[1014]= 32'b11111111111111111111111101011100;
    assign rom[1015]= 32'b11111111111111111111111101011011;
    assign rom[1016]= 32'b11111111111111111111111101011010;
    assign rom[1017]= 32'b11111111111111111111111101011001;
    assign rom[1018]= 32'b11111111111111111111111101011000;
    assign rom[1019]= 32'b11111111111111111111111101010111;
    assign rom[1020]= 32'b11111111111111111111111101010101;
    assign rom[1021]= 32'b11111111111111111111111101010100;
    assign rom[1022]= 32'b11111111111111111111111101010011;
    assign rom[1023]= 32'b11111111111111111111111101010010;
    assign rom[1024]= 32'b11111111111111111111111101010001;
    assign rom[1025]= 32'b11111111111111111111111101001111;
    assign rom[1026]= 32'b11111111111111111111111101001110;
    assign rom[1027]= 32'b11111111111111111111111101001101;
    assign rom[1028]= 32'b11111111111111111111111101001100;
    assign rom[1029]= 32'b11111111111111111111111101001011;
    assign rom[1030]= 32'b11111111111111111111111101001001;
    assign rom[1031]= 32'b11111111111111111111111101001000;
    assign rom[1032]= 32'b11111111111111111111111101000111;
    assign rom[1033]= 32'b11111111111111111111111101000110;
    assign rom[1034]= 32'b11111111111111111111111101000100;
    assign rom[1035]= 32'b11111111111111111111111101000011;
    assign rom[1036]= 32'b11111111111111111111111101000010;
    assign rom[1037]= 32'b11111111111111111111111101000000;
    assign rom[1038]= 32'b11111111111111111111111100111111;
    assign rom[1039]= 32'b11111111111111111111111100111110;
    assign rom[1040]= 32'b11111111111111111111111100111100;
    assign rom[1041]= 32'b11111111111111111111111100111011;
    assign rom[1042]= 32'b11111111111111111111111100111010;
    assign rom[1043]= 32'b11111111111111111111111100111000;
    assign rom[1044]= 32'b11111111111111111111111100110111;
    assign rom[1045]= 32'b11111111111111111111111100110110;
    assign rom[1046]= 32'b11111111111111111111111100110100;
    assign rom[1047]= 32'b11111111111111111111111100110011;
    assign rom[1048]= 32'b11111111111111111111111100110001;
    assign rom[1049]= 32'b11111111111111111111111100110000;
    assign rom[1050]= 32'b11111111111111111111111100101111;
    assign rom[1051]= 32'b11111111111111111111111100101101;
    assign rom[1052]= 32'b11111111111111111111111100101100;
    assign rom[1053]= 32'b11111111111111111111111100101010;
    assign rom[1054]= 32'b11111111111111111111111100101001;
    assign rom[1055]= 32'b11111111111111111111111100100111;
    assign rom[1056]= 32'b11111111111111111111111100100110;
    assign rom[1057]= 32'b11111111111111111111111100100100;
    assign rom[1058]= 32'b11111111111111111111111100100011;
    assign rom[1059]= 32'b11111111111111111111111100100001;
    assign rom[1060]= 32'b11111111111111111111111100100000;
    assign rom[1061]= 32'b11111111111111111111111100011110;
    assign rom[1062]= 32'b11111111111111111111111100011101;
    assign rom[1063]= 32'b11111111111111111111111100011011;
    assign rom[1064]= 32'b11111111111111111111111100011010;
    assign rom[1065]= 32'b11111111111111111111111100011000;
    assign rom[1066]= 32'b11111111111111111111111100010110;
    assign rom[1067]= 32'b11111111111111111111111100010101;
    assign rom[1068]= 32'b11111111111111111111111100010011;
    assign rom[1069]= 32'b11111111111111111111111100010010;
    assign rom[1070]= 32'b11111111111111111111111100010000;
    assign rom[1071]= 32'b11111111111111111111111100001110;
    assign rom[1072]= 32'b11111111111111111111111100001101;
    assign rom[1073]= 32'b11111111111111111111111100001011;
    assign rom[1074]= 32'b11111111111111111111111100001001;
    assign rom[1075]= 32'b11111111111111111111111100001000;
    assign rom[1076]= 32'b11111111111111111111111100000110;
    assign rom[1077]= 32'b11111111111111111111111100000100;
    assign rom[1078]= 32'b11111111111111111111111100000011;
    assign rom[1079]= 32'b11111111111111111111111100000001;
    assign rom[1080]= 32'b11111111111111111111111011111111;
    assign rom[1081]= 32'b11111111111111111111111011111101;
    assign rom[1082]= 32'b11111111111111111111111011111100;
    assign rom[1083]= 32'b11111111111111111111111011111010;
    assign rom[1084]= 32'b11111111111111111111111011111000;
    assign rom[1085]= 32'b11111111111111111111111011110110;
    assign rom[1086]= 32'b11111111111111111111111011110100;
    assign rom[1087]= 32'b11111111111111111111111011110011;
    assign rom[1088]= 32'b11111111111111111111111011110001;
    assign rom[1089]= 32'b11111111111111111111111011101111;
    assign rom[1090]= 32'b11111111111111111111111011101101;
    assign rom[1091]= 32'b11111111111111111111111011101011;
    assign rom[1092]= 32'b11111111111111111111111011101001;
    assign rom[1093]= 32'b11111111111111111111111011100111;
    assign rom[1094]= 32'b11111111111111111111111011100101;
    assign rom[1095]= 32'b11111111111111111111111011100100;
    assign rom[1096]= 32'b11111111111111111111111011100010;
    assign rom[1097]= 32'b11111111111111111111111011100000;
    assign rom[1098]= 32'b11111111111111111111111011011110;
    assign rom[1099]= 32'b11111111111111111111111011011100;
    assign rom[1100]= 32'b11111111111111111111111011011010;
    assign rom[1101]= 32'b11111111111111111111111011011000;
    assign rom[1102]= 32'b11111111111111111111111011010110;
    assign rom[1103]= 32'b11111111111111111111111011010100;
    assign rom[1104]= 32'b11111111111111111111111011010010;
    assign rom[1105]= 32'b11111111111111111111111011010000;
    assign rom[1106]= 32'b11111111111111111111111011001110;
    assign rom[1107]= 32'b11111111111111111111111011001011;
    assign rom[1108]= 32'b11111111111111111111111011001001;
    assign rom[1109]= 32'b11111111111111111111111011000111;
    assign rom[1110]= 32'b11111111111111111111111011000101;
    assign rom[1111]= 32'b11111111111111111111111011000011;
    assign rom[1112]= 32'b11111111111111111111111011000001;
    assign rom[1113]= 32'b11111111111111111111111010111111;
    assign rom[1114]= 32'b11111111111111111111111010111101;
    assign rom[1115]= 32'b11111111111111111111111010111010;
    assign rom[1116]= 32'b11111111111111111111111010111000;
    assign rom[1117]= 32'b11111111111111111111111010110110;
    assign rom[1118]= 32'b11111111111111111111111010110100;
    assign rom[1119]= 32'b11111111111111111111111010110001;
    assign rom[1120]= 32'b11111111111111111111111010101111;
    assign rom[1121]= 32'b11111111111111111111111010101101;
    assign rom[1122]= 32'b11111111111111111111111010101011;
    assign rom[1123]= 32'b11111111111111111111111010101000;
    assign rom[1124]= 32'b11111111111111111111111010100110;
    assign rom[1125]= 32'b11111111111111111111111010100100;
    assign rom[1126]= 32'b11111111111111111111111010100001;
    assign rom[1127]= 32'b11111111111111111111111010011111;
    assign rom[1128]= 32'b11111111111111111111111010011101;
    assign rom[1129]= 32'b11111111111111111111111010011010;
    assign rom[1130]= 32'b11111111111111111111111010011000;
    assign rom[1131]= 32'b11111111111111111111111010010101;
    assign rom[1132]= 32'b11111111111111111111111010010011;
    assign rom[1133]= 32'b11111111111111111111111010010000;
    assign rom[1134]= 32'b11111111111111111111111010001110;
    assign rom[1135]= 32'b11111111111111111111111010001011;
    assign rom[1136]= 32'b11111111111111111111111010001001;
    assign rom[1137]= 32'b11111111111111111111111010000110;
    assign rom[1138]= 32'b11111111111111111111111010000100;
    assign rom[1139]= 32'b11111111111111111111111010000001;
    assign rom[1140]= 32'b11111111111111111111111001111111;
    assign rom[1141]= 32'b11111111111111111111111001111100;
    assign rom[1142]= 32'b11111111111111111111111001111001;
    assign rom[1143]= 32'b11111111111111111111111001110111;
    assign rom[1144]= 32'b11111111111111111111111001110100;
    assign rom[1145]= 32'b11111111111111111111111001110010;
    assign rom[1146]= 32'b11111111111111111111111001101111;
    assign rom[1147]= 32'b11111111111111111111111001101100;
    assign rom[1148]= 32'b11111111111111111111111001101001;
    assign rom[1149]= 32'b11111111111111111111111001100111;
    assign rom[1150]= 32'b11111111111111111111111001100100;
    assign rom[1151]= 32'b11111111111111111111111001100001;
    assign rom[1152]= 32'b11111111111111111111111001011110;
    assign rom[1153]= 32'b11111111111111111111111001011100;
    assign rom[1154]= 32'b11111111111111111111111001011001;
    assign rom[1155]= 32'b11111111111111111111111001010110;
    assign rom[1156]= 32'b11111111111111111111111001010011;
    assign rom[1157]= 32'b11111111111111111111111001010000;
    assign rom[1158]= 32'b11111111111111111111111001001101;
    assign rom[1159]= 32'b11111111111111111111111001001010;
    assign rom[1160]= 32'b11111111111111111111111001000111;
    assign rom[1161]= 32'b11111111111111111111111001000100;
    assign rom[1162]= 32'b11111111111111111111111001000001;
    assign rom[1163]= 32'b11111111111111111111111000111110;
    assign rom[1164]= 32'b11111111111111111111111000111011;
    assign rom[1165]= 32'b11111111111111111111111000111000;
    assign rom[1166]= 32'b11111111111111111111111000110101;
    assign rom[1167]= 32'b11111111111111111111111000110010;
    assign rom[1168]= 32'b11111111111111111111111000101111;
    assign rom[1169]= 32'b11111111111111111111111000101100;
    assign rom[1170]= 32'b11111111111111111111111000101001;
    assign rom[1171]= 32'b11111111111111111111111000100110;
    assign rom[1172]= 32'b11111111111111111111111000100011;
    assign rom[1173]= 32'b11111111111111111111111000011111;
    assign rom[1174]= 32'b11111111111111111111111000011100;
    assign rom[1175]= 32'b11111111111111111111111000011001;
    assign rom[1176]= 32'b11111111111111111111111000010110;
    assign rom[1177]= 32'b11111111111111111111111000010010;
    assign rom[1178]= 32'b11111111111111111111111000001111;
    assign rom[1179]= 32'b11111111111111111111111000001100;
    assign rom[1180]= 32'b11111111111111111111111000001000;
    assign rom[1181]= 32'b11111111111111111111111000000101;
    assign rom[1182]= 32'b11111111111111111111111000000010;
    assign rom[1183]= 32'b11111111111111111111110111111110;
    assign rom[1184]= 32'b11111111111111111111110111111011;
    assign rom[1185]= 32'b11111111111111111111110111110111;
    assign rom[1186]= 32'b11111111111111111111110111110100;
    assign rom[1187]= 32'b11111111111111111111110111110000;
    assign rom[1188]= 32'b11111111111111111111110111101101;
    assign rom[1189]= 32'b11111111111111111111110111101001;
    assign rom[1190]= 32'b11111111111111111111110111100110;
    assign rom[1191]= 32'b11111111111111111111110111100010;
    assign rom[1192]= 32'b11111111111111111111110111011111;
    assign rom[1193]= 32'b11111111111111111111110111011011;
    assign rom[1194]= 32'b11111111111111111111110111010111;
    assign rom[1195]= 32'b11111111111111111111110111010100;
    assign rom[1196]= 32'b11111111111111111111110111010000;
    assign rom[1197]= 32'b11111111111111111111110111001100;
    assign rom[1198]= 32'b11111111111111111111110111001000;
    assign rom[1199]= 32'b11111111111111111111110111000101;
    assign rom[1200]= 32'b11111111111111111111110111000001;
    assign rom[1201]= 32'b11111111111111111111110110111101;
    assign rom[1202]= 32'b11111111111111111111110110111001;
    assign rom[1203]= 32'b11111111111111111111110110110101;
    assign rom[1204]= 32'b11111111111111111111110110110001;
    assign rom[1205]= 32'b11111111111111111111110110101101;
    assign rom[1206]= 32'b11111111111111111111110110101001;
    assign rom[1207]= 32'b11111111111111111111110110100110;
    assign rom[1208]= 32'b11111111111111111111110110100010;
    assign rom[1209]= 32'b11111111111111111111110110011101;
    assign rom[1210]= 32'b11111111111111111111110110011001;
    assign rom[1211]= 32'b11111111111111111111110110010101;
    assign rom[1212]= 32'b11111111111111111111110110010001;
    assign rom[1213]= 32'b11111111111111111111110110001101;
    assign rom[1214]= 32'b11111111111111111111110110001001;
    assign rom[1215]= 32'b11111111111111111111110110000101;
    assign rom[1216]= 32'b11111111111111111111110110000001;
    assign rom[1217]= 32'b11111111111111111111110101111100;
    assign rom[1218]= 32'b11111111111111111111110101111000;
    assign rom[1219]= 32'b11111111111111111111110101110100;
    assign rom[1220]= 32'b11111111111111111111110101101111;
    assign rom[1221]= 32'b11111111111111111111110101101011;
    assign rom[1222]= 32'b11111111111111111111110101100111;
    assign rom[1223]= 32'b11111111111111111111110101100010;
    assign rom[1224]= 32'b11111111111111111111110101011110;
    assign rom[1225]= 32'b11111111111111111111110101011001;
    assign rom[1226]= 32'b11111111111111111111110101010101;
    assign rom[1227]= 32'b11111111111111111111110101010000;
    assign rom[1228]= 32'b11111111111111111111110101001100;
    assign rom[1229]= 32'b11111111111111111111110101000111;
    assign rom[1230]= 32'b11111111111111111111110101000011;
    assign rom[1231]= 32'b11111111111111111111110100111110;
    assign rom[1232]= 32'b11111111111111111111110100111001;
    assign rom[1233]= 32'b11111111111111111111110100110101;
    assign rom[1234]= 32'b11111111111111111111110100110000;
    assign rom[1235]= 32'b11111111111111111111110100101011;
    assign rom[1236]= 32'b11111111111111111111110100100110;
    assign rom[1237]= 32'b11111111111111111111110100100010;
    assign rom[1238]= 32'b11111111111111111111110100011101;
    assign rom[1239]= 32'b11111111111111111111110100011000;
    assign rom[1240]= 32'b11111111111111111111110100010011;
    assign rom[1241]= 32'b11111111111111111111110100001110;
    assign rom[1242]= 32'b11111111111111111111110100001001;
    assign rom[1243]= 32'b11111111111111111111110100000100;
    assign rom[1244]= 32'b11111111111111111111110011111111;
    assign rom[1245]= 32'b11111111111111111111110011111010;
    assign rom[1246]= 32'b11111111111111111111110011110101;
    assign rom[1247]= 32'b11111111111111111111110011110000;
    assign rom[1248]= 32'b11111111111111111111110011101011;
    assign rom[1249]= 32'b11111111111111111111110011100101;
    assign rom[1250]= 32'b11111111111111111111110011100000;
    assign rom[1251]= 32'b11111111111111111111110011011011;
    assign rom[1252]= 32'b11111111111111111111110011010110;
    assign rom[1253]= 32'b11111111111111111111110011010000;
    assign rom[1254]= 32'b11111111111111111111110011001011;
    assign rom[1255]= 32'b11111111111111111111110011000101;
    assign rom[1256]= 32'b11111111111111111111110011000000;
    assign rom[1257]= 32'b11111111111111111111110010111011;
    assign rom[1258]= 32'b11111111111111111111110010110101;
    assign rom[1259]= 32'b11111111111111111111110010110000;
    assign rom[1260]= 32'b11111111111111111111110010101010;
    assign rom[1261]= 32'b11111111111111111111110010100100;
    assign rom[1262]= 32'b11111111111111111111110010011111;
    assign rom[1263]= 32'b11111111111111111111110010011001;
    assign rom[1264]= 32'b11111111111111111111110010010011;
    assign rom[1265]= 32'b11111111111111111111110010001110;
    assign rom[1266]= 32'b11111111111111111111110010001000;
    assign rom[1267]= 32'b11111111111111111111110010000010;
    assign rom[1268]= 32'b11111111111111111111110001111100;
    assign rom[1269]= 32'b11111111111111111111110001110110;
    assign rom[1270]= 32'b11111111111111111111110001110000;
    assign rom[1271]= 32'b11111111111111111111110001101010;
    assign rom[1272]= 32'b11111111111111111111110001100100;
    assign rom[1273]= 32'b11111111111111111111110001011110;
    assign rom[1274]= 32'b11111111111111111111110001011000;
    assign rom[1275]= 32'b11111111111111111111110001010010;
    assign rom[1276]= 32'b11111111111111111111110001001100;
    assign rom[1277]= 32'b11111111111111111111110001000110;
    assign rom[1278]= 32'b11111111111111111111110001000000;
    assign rom[1279]= 32'b11111111111111111111110000111001;
    assign rom[1280]= 32'b11111111111111111111110000110011;
    assign rom[1281]= 32'b11111111111111111111110000101101;
    assign rom[1282]= 32'b11111111111111111111110000100110;
    assign rom[1283]= 32'b11111111111111111111110000100000;
    assign rom[1284]= 32'b11111111111111111111110000011001;
    assign rom[1285]= 32'b11111111111111111111110000010011;
    assign rom[1286]= 32'b11111111111111111111110000001100;
    assign rom[1287]= 32'b11111111111111111111110000000110;
    assign rom[1288]= 32'b11111111111111111111101111111111;
    assign rom[1289]= 32'b11111111111111111111101111111000;
    assign rom[1290]= 32'b11111111111111111111101111110010;
    assign rom[1291]= 32'b11111111111111111111101111101011;
    assign rom[1292]= 32'b11111111111111111111101111100100;
    assign rom[1293]= 32'b11111111111111111111101111011101;
    assign rom[1294]= 32'b11111111111111111111101111010110;
    assign rom[1295]= 32'b11111111111111111111101111010000;
    assign rom[1296]= 32'b11111111111111111111101111001001;
    assign rom[1297]= 32'b11111111111111111111101111000010;
    assign rom[1298]= 32'b11111111111111111111101110111011;
    assign rom[1299]= 32'b11111111111111111111101110110011;
    assign rom[1300]= 32'b11111111111111111111101110101100;
    assign rom[1301]= 32'b11111111111111111111101110100101;
    assign rom[1302]= 32'b11111111111111111111101110011110;
    assign rom[1303]= 32'b11111111111111111111101110010111;
    assign rom[1304]= 32'b11111111111111111111101110001111;
    assign rom[1305]= 32'b11111111111111111111101110001000;
    assign rom[1306]= 32'b11111111111111111111101110000000;
    assign rom[1307]= 32'b11111111111111111111101101111001;
    assign rom[1308]= 32'b11111111111111111111101101110010;
    assign rom[1309]= 32'b11111111111111111111101101101010;
    assign rom[1310]= 32'b11111111111111111111101101100010;
    assign rom[1311]= 32'b11111111111111111111101101011011;
    assign rom[1312]= 32'b11111111111111111111101101010011;
    assign rom[1313]= 32'b11111111111111111111101101001011;
    assign rom[1314]= 32'b11111111111111111111101101000100;
    assign rom[1315]= 32'b11111111111111111111101100111100;
    assign rom[1316]= 32'b11111111111111111111101100110100;
    assign rom[1317]= 32'b11111111111111111111101100101100;
    assign rom[1318]= 32'b11111111111111111111101100100100;
    assign rom[1319]= 32'b11111111111111111111101100011100;
    assign rom[1320]= 32'b11111111111111111111101100010100;
    assign rom[1321]= 32'b11111111111111111111101100001100;
    assign rom[1322]= 32'b11111111111111111111101100000011;
    assign rom[1323]= 32'b11111111111111111111101011111011;
    assign rom[1324]= 32'b11111111111111111111101011110011;
    assign rom[1325]= 32'b11111111111111111111101011101011;
    assign rom[1326]= 32'b11111111111111111111101011100010;
    assign rom[1327]= 32'b11111111111111111111101011011010;
    assign rom[1328]= 32'b11111111111111111111101011010001;
    assign rom[1329]= 32'b11111111111111111111101011001001;
    assign rom[1330]= 32'b11111111111111111111101011000000;
    assign rom[1331]= 32'b11111111111111111111101010111000;
    assign rom[1332]= 32'b11111111111111111111101010101111;
    assign rom[1333]= 32'b11111111111111111111101010100110;
    assign rom[1334]= 32'b11111111111111111111101010011101;
    assign rom[1335]= 32'b11111111111111111111101010010101;
    assign rom[1336]= 32'b11111111111111111111101010001100;
    assign rom[1337]= 32'b11111111111111111111101010000011;
    assign rom[1338]= 32'b11111111111111111111101001111010;
    assign rom[1339]= 32'b11111111111111111111101001110001;
    assign rom[1340]= 32'b11111111111111111111101001100111;
    assign rom[1341]= 32'b11111111111111111111101001011110;
    assign rom[1342]= 32'b11111111111111111111101001010101;
    assign rom[1343]= 32'b11111111111111111111101001001100;
    assign rom[1344]= 32'b11111111111111111111101001000010;
    assign rom[1345]= 32'b11111111111111111111101000111001;
    assign rom[1346]= 32'b11111111111111111111101000110000;
    assign rom[1347]= 32'b11111111111111111111101000100110;
    assign rom[1348]= 32'b11111111111111111111101000011100;
    assign rom[1349]= 32'b11111111111111111111101000010011;
    assign rom[1350]= 32'b11111111111111111111101000001001;
    assign rom[1351]= 32'b11111111111111111111100111111111;
    assign rom[1352]= 32'b11111111111111111111100111110110;
    assign rom[1353]= 32'b11111111111111111111100111101100;
    assign rom[1354]= 32'b11111111111111111111100111100010;
    assign rom[1355]= 32'b11111111111111111111100111011000;
    assign rom[1356]= 32'b11111111111111111111100111001110;
    assign rom[1357]= 32'b11111111111111111111100111000100;
    assign rom[1358]= 32'b11111111111111111111100110111010;
    assign rom[1359]= 32'b11111111111111111111100110101111;
    assign rom[1360]= 32'b11111111111111111111100110100101;
    assign rom[1361]= 32'b11111111111111111111100110011011;
    assign rom[1362]= 32'b11111111111111111111100110010000;
    assign rom[1363]= 32'b11111111111111111111100110000110;
    assign rom[1364]= 32'b11111111111111111111100101111011;
    assign rom[1365]= 32'b11111111111111111111100101110001;
    assign rom[1366]= 32'b11111111111111111111100101100110;
    assign rom[1367]= 32'b11111111111111111111100101011011;
    assign rom[1368]= 32'b11111111111111111111100101010000;
    assign rom[1369]= 32'b11111111111111111111100101000110;
    assign rom[1370]= 32'b11111111111111111111100100111011;
    assign rom[1371]= 32'b11111111111111111111100100110000;
    assign rom[1372]= 32'b11111111111111111111100100100101;
    assign rom[1373]= 32'b11111111111111111111100100011010;
    assign rom[1374]= 32'b11111111111111111111100100001110;
    assign rom[1375]= 32'b11111111111111111111100100000011;
    assign rom[1376]= 32'b11111111111111111111100011111000;
    assign rom[1377]= 32'b11111111111111111111100011101100;
    assign rom[1378]= 32'b11111111111111111111100011100001;
    assign rom[1379]= 32'b11111111111111111111100011010101;
    assign rom[1380]= 32'b11111111111111111111100011001010;
    assign rom[1381]= 32'b11111111111111111111100010111110;
    assign rom[1382]= 32'b11111111111111111111100010110010;
    assign rom[1383]= 32'b11111111111111111111100010100111;
    assign rom[1384]= 32'b11111111111111111111100010011011;
    assign rom[1385]= 32'b11111111111111111111100010001111;
    assign rom[1386]= 32'b11111111111111111111100010000011;
    assign rom[1387]= 32'b11111111111111111111100001110111;
    assign rom[1388]= 32'b11111111111111111111100001101011;
    assign rom[1389]= 32'b11111111111111111111100001011110;
    assign rom[1390]= 32'b11111111111111111111100001010010;
    assign rom[1391]= 32'b11111111111111111111100001000110;
    assign rom[1392]= 32'b11111111111111111111100000111001;
    assign rom[1393]= 32'b11111111111111111111100000101101;
    assign rom[1394]= 32'b11111111111111111111100000100000;
    assign rom[1395]= 32'b11111111111111111111100000010100;
    assign rom[1396]= 32'b11111111111111111111100000000111;
    assign rom[1397]= 32'b11111111111111111111011111111010;
    assign rom[1398]= 32'b11111111111111111111011111101101;
    assign rom[1399]= 32'b11111111111111111111011111100000;
    assign rom[1400]= 32'b11111111111111111111011111010011;
    assign rom[1401]= 32'b11111111111111111111011111000110;
    assign rom[1402]= 32'b11111111111111111111011110111001;
    assign rom[1403]= 32'b11111111111111111111011110101100;
    assign rom[1404]= 32'b11111111111111111111011110011110;
    assign rom[1405]= 32'b11111111111111111111011110010001;
    assign rom[1406]= 32'b11111111111111111111011110000011;
    assign rom[1407]= 32'b11111111111111111111011101110110;
    assign rom[1408]= 32'b11111111111111111111011101101000;
    assign rom[1409]= 32'b11111111111111111111011101011010;
    assign rom[1410]= 32'b11111111111111111111011101001100;
    assign rom[1411]= 32'b11111111111111111111011100111111;
    assign rom[1412]= 32'b11111111111111111111011100110001;
    assign rom[1413]= 32'b11111111111111111111011100100011;
    assign rom[1414]= 32'b11111111111111111111011100010100;
    assign rom[1415]= 32'b11111111111111111111011100000110;
    assign rom[1416]= 32'b11111111111111111111011011111000;
    assign rom[1417]= 32'b11111111111111111111011011101010;
    assign rom[1418]= 32'b11111111111111111111011011011011;
    assign rom[1419]= 32'b11111111111111111111011011001101;
    assign rom[1420]= 32'b11111111111111111111011010111110;
    assign rom[1421]= 32'b11111111111111111111011010101111;
    assign rom[1422]= 32'b11111111111111111111011010100000;
    assign rom[1423]= 32'b11111111111111111111011010010001;
    assign rom[1424]= 32'b11111111111111111111011010000010;
    assign rom[1425]= 32'b11111111111111111111011001110011;
    assign rom[1426]= 32'b11111111111111111111011001100100;
    assign rom[1427]= 32'b11111111111111111111011001010101;
    assign rom[1428]= 32'b11111111111111111111011001000110;
    assign rom[1429]= 32'b11111111111111111111011000110110;
    assign rom[1430]= 32'b11111111111111111111011000100111;
    assign rom[1431]= 32'b11111111111111111111011000010111;
    assign rom[1432]= 32'b11111111111111111111011000001000;
    assign rom[1433]= 32'b11111111111111111111010111111000;
    assign rom[1434]= 32'b11111111111111111111010111101000;
    assign rom[1435]= 32'b11111111111111111111010111011000;
    assign rom[1436]= 32'b11111111111111111111010111001000;
    assign rom[1437]= 32'b11111111111111111111010110111000;
    assign rom[1438]= 32'b11111111111111111111010110101000;
    assign rom[1439]= 32'b11111111111111111111010110010111;
    assign rom[1440]= 32'b11111111111111111111010110000111;
    assign rom[1441]= 32'b11111111111111111111010101110110;
    assign rom[1442]= 32'b11111111111111111111010101100110;
    assign rom[1443]= 32'b11111111111111111111010101010101;
    assign rom[1444]= 32'b11111111111111111111010101000100;
    assign rom[1445]= 32'b11111111111111111111010100110011;
    assign rom[1446]= 32'b11111111111111111111010100100011;
    assign rom[1447]= 32'b11111111111111111111010100010001;
    assign rom[1448]= 32'b11111111111111111111010100000000;
    assign rom[1449]= 32'b11111111111111111111010011101111;
    assign rom[1450]= 32'b11111111111111111111010011011110;
    assign rom[1451]= 32'b11111111111111111111010011001100;
    assign rom[1452]= 32'b11111111111111111111010010111011;
    assign rom[1453]= 32'b11111111111111111111010010101001;
    assign rom[1454]= 32'b11111111111111111111010010010111;
    assign rom[1455]= 32'b11111111111111111111010010000101;
    assign rom[1456]= 32'b11111111111111111111010001110100;
    assign rom[1457]= 32'b11111111111111111111010001100001;
    assign rom[1458]= 32'b11111111111111111111010001001111;
    assign rom[1459]= 32'b11111111111111111111010000111101;
    assign rom[1460]= 32'b11111111111111111111010000101011;
    assign rom[1461]= 32'b11111111111111111111010000011000;
    assign rom[1462]= 32'b11111111111111111111010000000110;
    assign rom[1463]= 32'b11111111111111111111001111110011;
    assign rom[1464]= 32'b11111111111111111111001111100000;
    assign rom[1465]= 32'b11111111111111111111001111001101;
    assign rom[1466]= 32'b11111111111111111111001110111011;
    assign rom[1467]= 32'b11111111111111111111001110100111;
    assign rom[1468]= 32'b11111111111111111111001110010100;
    assign rom[1469]= 32'b11111111111111111111001110000001;
    assign rom[1470]= 32'b11111111111111111111001101101110;
    assign rom[1471]= 32'b11111111111111111111001101011010;
    assign rom[1472]= 32'b11111111111111111111001101000111;
    assign rom[1473]= 32'b11111111111111111111001100110011;
    assign rom[1474]= 32'b11111111111111111111001100011111;
    assign rom[1475]= 32'b11111111111111111111001100001011;
    assign rom[1476]= 32'b11111111111111111111001011110111;
    assign rom[1477]= 32'b11111111111111111111001011100011;
    assign rom[1478]= 32'b11111111111111111111001011001111;
    assign rom[1479]= 32'b11111111111111111111001010111010;
    assign rom[1480]= 32'b11111111111111111111001010100110;
    assign rom[1481]= 32'b11111111111111111111001010010001;
    assign rom[1482]= 32'b11111111111111111111001001111101;
    assign rom[1483]= 32'b11111111111111111111001001101000;
    assign rom[1484]= 32'b11111111111111111111001001010011;
    assign rom[1485]= 32'b11111111111111111111001000111110;
    assign rom[1486]= 32'b11111111111111111111001000101001;
    assign rom[1487]= 32'b11111111111111111111001000010011;
    assign rom[1488]= 32'b11111111111111111111000111111110;
    assign rom[1489]= 32'b11111111111111111111000111101000;
    assign rom[1490]= 32'b11111111111111111111000111010011;
    assign rom[1491]= 32'b11111111111111111111000110111101;
    assign rom[1492]= 32'b11111111111111111111000110100111;
    assign rom[1493]= 32'b11111111111111111111000110010001;
    assign rom[1494]= 32'b11111111111111111111000101111011;
    assign rom[1495]= 32'b11111111111111111111000101100101;
    assign rom[1496]= 32'b11111111111111111111000101001111;
    assign rom[1497]= 32'b11111111111111111111000100111000;
    assign rom[1498]= 32'b11111111111111111111000100100010;
    assign rom[1499]= 32'b11111111111111111111000100001011;
    assign rom[1500]= 32'b11111111111111111111000011110100;
    assign rom[1501]= 32'b11111111111111111111000011011101;
    assign rom[1502]= 32'b11111111111111111111000011000110;
    assign rom[1503]= 32'b11111111111111111111000010101111;
    assign rom[1504]= 32'b11111111111111111111000010011000;
    assign rom[1505]= 32'b11111111111111111111000010000000;
    assign rom[1506]= 32'b11111111111111111111000001101001;
    assign rom[1507]= 32'b11111111111111111111000001010001;
    assign rom[1508]= 32'b11111111111111111111000000111001;
    assign rom[1509]= 32'b11111111111111111111000000100010;
    assign rom[1510]= 32'b11111111111111111111000000001010;
    assign rom[1511]= 32'b11111111111111111110111111110001;
    assign rom[1512]= 32'b11111111111111111110111111011001;
    assign rom[1513]= 32'b11111111111111111110111111000001;
    assign rom[1514]= 32'b11111111111111111110111110101000;
    assign rom[1515]= 32'b11111111111111111110111110001111;
    assign rom[1516]= 32'b11111111111111111110111101110111;
    assign rom[1517]= 32'b11111111111111111110111101011110;
    assign rom[1518]= 32'b11111111111111111110111101000101;
    assign rom[1519]= 32'b11111111111111111110111100101100;
    assign rom[1520]= 32'b11111111111111111110111100010010;
    assign rom[1521]= 32'b11111111111111111110111011111001;
    assign rom[1522]= 32'b11111111111111111110111011011111;
    assign rom[1523]= 32'b11111111111111111110111011000110;
    assign rom[1524]= 32'b11111111111111111110111010101100;
    assign rom[1525]= 32'b11111111111111111110111010010010;
    assign rom[1526]= 32'b11111111111111111110111001111000;
    assign rom[1527]= 32'b11111111111111111110111001011101;
    assign rom[1528]= 32'b11111111111111111110111001000011;
    assign rom[1529]= 32'b11111111111111111110111000101000;
    assign rom[1530]= 32'b11111111111111111110111000001110;
    assign rom[1531]= 32'b11111111111111111110110111110011;
    assign rom[1532]= 32'b11111111111111111110110111011000;
    assign rom[1533]= 32'b11111111111111111110110110111101;
    assign rom[1534]= 32'b11111111111111111110110110100010;
    assign rom[1535]= 32'b11111111111111111110110110000111;
    assign rom[1536]= 32'b11111111111111111110110101101011;
    assign rom[1537]= 32'b11111111111111111110110101010000;
    assign rom[1538]= 32'b11111111111111111110110100110100;
    assign rom[1539]= 32'b11111111111111111110110100011000;
    assign rom[1540]= 32'b11111111111111111110110011111100;
    assign rom[1541]= 32'b11111111111111111110110011100000;
    assign rom[1542]= 32'b11111111111111111110110011000011;
    assign rom[1543]= 32'b11111111111111111110110010100111;
    assign rom[1544]= 32'b11111111111111111110110010001010;
    assign rom[1545]= 32'b11111111111111111110110001101110;
    assign rom[1546]= 32'b11111111111111111110110001010001;
    assign rom[1547]= 32'b11111111111111111110110000110100;
    assign rom[1548]= 32'b11111111111111111110110000010111;
    assign rom[1549]= 32'b11111111111111111110101111111001;
    assign rom[1550]= 32'b11111111111111111110101111011100;
    assign rom[1551]= 32'b11111111111111111110101110111110;
    assign rom[1552]= 32'b11111111111111111110101110100001;
    assign rom[1553]= 32'b11111111111111111110101110000011;
    assign rom[1554]= 32'b11111111111111111110101101100101;
    assign rom[1555]= 32'b11111111111111111110101101000110;
    assign rom[1556]= 32'b11111111111111111110101100101000;
    assign rom[1557]= 32'b11111111111111111110101100001010;
    assign rom[1558]= 32'b11111111111111111110101011101011;
    assign rom[1559]= 32'b11111111111111111110101011001100;
    assign rom[1560]= 32'b11111111111111111110101010101101;
    assign rom[1561]= 32'b11111111111111111110101010001110;
    assign rom[1562]= 32'b11111111111111111110101001101111;
    assign rom[1563]= 32'b11111111111111111110101001010000;
    assign rom[1564]= 32'b11111111111111111110101000110000;
    assign rom[1565]= 32'b11111111111111111110101000010001;
    assign rom[1566]= 32'b11111111111111111110100111110001;
    assign rom[1567]= 32'b11111111111111111110100111010001;
    assign rom[1568]= 32'b11111111111111111110100110110001;
    assign rom[1569]= 32'b11111111111111111110100110010000;
    assign rom[1570]= 32'b11111111111111111110100101110000;
    assign rom[1571]= 32'b11111111111111111110100101001111;
    assign rom[1572]= 32'b11111111111111111110100100101111;
    assign rom[1573]= 32'b11111111111111111110100100001110;
    assign rom[1574]= 32'b11111111111111111110100011101101;
    assign rom[1575]= 32'b11111111111111111110100011001100;
    assign rom[1576]= 32'b11111111111111111110100010101010;
    assign rom[1577]= 32'b11111111111111111110100010001001;
    assign rom[1578]= 32'b11111111111111111110100001100111;
    assign rom[1579]= 32'b11111111111111111110100001000101;
    assign rom[1580]= 32'b11111111111111111110100000100011;
    assign rom[1581]= 32'b11111111111111111110100000000001;
    assign rom[1582]= 32'b11111111111111111110011111011111;
    assign rom[1583]= 32'b11111111111111111110011110111100;
    assign rom[1584]= 32'b11111111111111111110011110011010;
    assign rom[1585]= 32'b11111111111111111110011101110111;
    assign rom[1586]= 32'b11111111111111111110011101010100;
    assign rom[1587]= 32'b11111111111111111110011100110001;
    assign rom[1588]= 32'b11111111111111111110011100001110;
    assign rom[1589]= 32'b11111111111111111110011011101010;
    assign rom[1590]= 32'b11111111111111111110011011000111;
    assign rom[1591]= 32'b11111111111111111110011010100011;
    assign rom[1592]= 32'b11111111111111111110011001111111;
    assign rom[1593]= 32'b11111111111111111110011001011011;
    assign rom[1594]= 32'b11111111111111111110011000110111;
    assign rom[1595]= 32'b11111111111111111110011000010011;
    assign rom[1596]= 32'b11111111111111111110010111101110;
    assign rom[1597]= 32'b11111111111111111110010111001010;
    assign rom[1598]= 32'b11111111111111111110010110100101;
    assign rom[1599]= 32'b11111111111111111110010110000000;
    assign rom[1600]= 32'b11111111111111111110010101011010;
    assign rom[1601]= 32'b11111111111111111110010100110101;
    assign rom[1602]= 32'b11111111111111111110010100010000;
    assign rom[1603]= 32'b11111111111111111110010011101010;
    assign rom[1604]= 32'b11111111111111111110010011000100;
    assign rom[1605]= 32'b11111111111111111110010010011110;
    assign rom[1606]= 32'b11111111111111111110010001111000;
    assign rom[1607]= 32'b11111111111111111110010001010010;
    assign rom[1608]= 32'b11111111111111111110010000101011;
    assign rom[1609]= 32'b11111111111111111110010000000101;
    assign rom[1610]= 32'b11111111111111111110001111011110;
    assign rom[1611]= 32'b11111111111111111110001110110111;
    assign rom[1612]= 32'b11111111111111111110001110010000;
    assign rom[1613]= 32'b11111111111111111110001101101000;
    assign rom[1614]= 32'b11111111111111111110001101000001;
    assign rom[1615]= 32'b11111111111111111110001100011001;
    assign rom[1616]= 32'b11111111111111111110001011110001;
    assign rom[1617]= 32'b11111111111111111110001011001001;
    assign rom[1618]= 32'b11111111111111111110001010100001;
    assign rom[1619]= 32'b11111111111111111110001001111001;
    assign rom[1620]= 32'b11111111111111111110001001010001;
    assign rom[1621]= 32'b11111111111111111110001000101000;
    assign rom[1622]= 32'b11111111111111111110000111111111;
    assign rom[1623]= 32'b11111111111111111110000111010110;
    assign rom[1624]= 32'b11111111111111111110000110101101;
    assign rom[1625]= 32'b11111111111111111110000110000100;
    assign rom[1626]= 32'b11111111111111111110000101011010;
    assign rom[1627]= 32'b11111111111111111110000100110001;
    assign rom[1628]= 32'b11111111111111111110000100000111;
    assign rom[1629]= 32'b11111111111111111110000011011101;
    assign rom[1630]= 32'b11111111111111111110000010110011;
    assign rom[1631]= 32'b11111111111111111110000010001000;
    assign rom[1632]= 32'b11111111111111111110000001011110;
    assign rom[1633]= 32'b11111111111111111110000000110011;
    assign rom[1634]= 32'b11111111111111111110000000001000;
    assign rom[1635]= 32'b11111111111111111101111111011101;
    assign rom[1636]= 32'b11111111111111111101111110110010;
    assign rom[1637]= 32'b11111111111111111101111110000111;
    assign rom[1638]= 32'b11111111111111111101111101011100;
    assign rom[1639]= 32'b11111111111111111101111100110000;
    assign rom[1640]= 32'b11111111111111111101111100000100;
    assign rom[1641]= 32'b11111111111111111101111011011000;
    assign rom[1642]= 32'b11111111111111111101111010101100;
    assign rom[1643]= 32'b11111111111111111101111010000000;
    assign rom[1644]= 32'b11111111111111111101111001010011;
    assign rom[1645]= 32'b11111111111111111101111000100111;
    assign rom[1646]= 32'b11111111111111111101110111111010;
    assign rom[1647]= 32'b11111111111111111101110111001101;
    assign rom[1648]= 32'b11111111111111111101110110100000;
    assign rom[1649]= 32'b11111111111111111101110101110010;
    assign rom[1650]= 32'b11111111111111111101110101000101;
    assign rom[1651]= 32'b11111111111111111101110100010111;
    assign rom[1652]= 32'b11111111111111111101110011101010;
    assign rom[1653]= 32'b11111111111111111101110010111100;
    assign rom[1654]= 32'b11111111111111111101110010001101;
    assign rom[1655]= 32'b11111111111111111101110001011111;
    assign rom[1656]= 32'b11111111111111111101110000110001;
    assign rom[1657]= 32'b11111111111111111101110000000010;
    assign rom[1658]= 32'b11111111111111111101101111010011;
    assign rom[1659]= 32'b11111111111111111101101110100100;
    assign rom[1660]= 32'b11111111111111111101101101110101;
    assign rom[1661]= 32'b11111111111111111101101101000110;
    assign rom[1662]= 32'b11111111111111111101101100010111;
    assign rom[1663]= 32'b11111111111111111101101011100111;
    assign rom[1664]= 32'b11111111111111111101101010110111;
    assign rom[1665]= 32'b11111111111111111101101010000111;
    assign rom[1666]= 32'b11111111111111111101101001010111;
    assign rom[1667]= 32'b11111111111111111101101000100111;
    assign rom[1668]= 32'b11111111111111111101100111110111;
    assign rom[1669]= 32'b11111111111111111101100111000110;
    assign rom[1670]= 32'b11111111111111111101100110010110;
    assign rom[1671]= 32'b11111111111111111101100101100101;
    assign rom[1672]= 32'b11111111111111111101100100110100;
    assign rom[1673]= 32'b11111111111111111101100100000011;
    assign rom[1674]= 32'b11111111111111111101100011010001;
    assign rom[1675]= 32'b11111111111111111101100010100000;
    assign rom[1676]= 32'b11111111111111111101100001101110;
    assign rom[1677]= 32'b11111111111111111101100000111100;
    assign rom[1678]= 32'b11111111111111111101100000001010;
    assign rom[1679]= 32'b11111111111111111101011111011000;
    assign rom[1680]= 32'b11111111111111111101011110100110;
    assign rom[1681]= 32'b11111111111111111101011101110100;
    assign rom[1682]= 32'b11111111111111111101011101000001;
    assign rom[1683]= 32'b11111111111111111101011100001111;
    assign rom[1684]= 32'b11111111111111111101011011011100;
    assign rom[1685]= 32'b11111111111111111101011010101001;
    assign rom[1686]= 32'b11111111111111111101011001110110;
    assign rom[1687]= 32'b11111111111111111101011001000010;
    assign rom[1688]= 32'b11111111111111111101011000001111;
    assign rom[1689]= 32'b11111111111111111101010111011011;
    assign rom[1690]= 32'b11111111111111111101010110101000;
    assign rom[1691]= 32'b11111111111111111101010101110100;
    assign rom[1692]= 32'b11111111111111111101010101000000;
    assign rom[1693]= 32'b11111111111111111101010100001100;
    assign rom[1694]= 32'b11111111111111111101010011011000;
    assign rom[1695]= 32'b11111111111111111101010010100011;
    assign rom[1696]= 32'b11111111111111111101010001101111;
    assign rom[1697]= 32'b11111111111111111101010000111010;
    assign rom[1698]= 32'b11111111111111111101010000000101;
    assign rom[1699]= 32'b11111111111111111101001111010000;
    assign rom[1700]= 32'b11111111111111111101001110011011;
    assign rom[1701]= 32'b11111111111111111101001101100110;
    assign rom[1702]= 32'b11111111111111111101001100110001;
    assign rom[1703]= 32'b11111111111111111101001011111011;
    assign rom[1704]= 32'b11111111111111111101001011000110;
    assign rom[1705]= 32'b11111111111111111101001010010000;
    assign rom[1706]= 32'b11111111111111111101001001011010;
    assign rom[1707]= 32'b11111111111111111101001000100100;
    assign rom[1708]= 32'b11111111111111111101000111101110;
    assign rom[1709]= 32'b11111111111111111101000110111000;
    assign rom[1710]= 32'b11111111111111111101000110000010;
    assign rom[1711]= 32'b11111111111111111101000101001011;
    assign rom[1712]= 32'b11111111111111111101000100010101;
    assign rom[1713]= 32'b11111111111111111101000011011110;
    assign rom[1714]= 32'b11111111111111111101000010100111;
    assign rom[1715]= 32'b11111111111111111101000001110001;
    assign rom[1716]= 32'b11111111111111111101000000111010;
    assign rom[1717]= 32'b11111111111111111101000000000010;
    assign rom[1718]= 32'b11111111111111111100111111001011;
    assign rom[1719]= 32'b11111111111111111100111110010100;
    assign rom[1720]= 32'b11111111111111111100111101011101;
    assign rom[1721]= 32'b11111111111111111100111100100101;
    assign rom[1722]= 32'b11111111111111111100111011101101;
    assign rom[1723]= 32'b11111111111111111100111010110110;
    assign rom[1724]= 32'b11111111111111111100111001111110;
    assign rom[1725]= 32'b11111111111111111100111001000110;
    assign rom[1726]= 32'b11111111111111111100111000001110;
    assign rom[1727]= 32'b11111111111111111100110111010110;
    assign rom[1728]= 32'b11111111111111111100110110011110;
    assign rom[1729]= 32'b11111111111111111100110101100110;
    assign rom[1730]= 32'b11111111111111111100110100101101;
    assign rom[1731]= 32'b11111111111111111100110011110101;
    assign rom[1732]= 32'b11111111111111111100110010111101;
    assign rom[1733]= 32'b11111111111111111100110010000100;
    assign rom[1734]= 32'b11111111111111111100110001001011;
    assign rom[1735]= 32'b11111111111111111100110000010011;
    assign rom[1736]= 32'b11111111111111111100101111011010;
    assign rom[1737]= 32'b11111111111111111100101110100001;
    assign rom[1738]= 32'b11111111111111111100101101101000;
    assign rom[1739]= 32'b11111111111111111100101100101111;
    assign rom[1740]= 32'b11111111111111111100101011110110;
    assign rom[1741]= 32'b11111111111111111100101010111101;
    assign rom[1742]= 32'b11111111111111111100101010000100;
    assign rom[1743]= 32'b11111111111111111100101001001011;
    assign rom[1744]= 32'b11111111111111111100101000010010;
    assign rom[1745]= 32'b11111111111111111100100111011000;
    assign rom[1746]= 32'b11111111111111111100100110011111;
    assign rom[1747]= 32'b11111111111111111100100101100110;
    assign rom[1748]= 32'b11111111111111111100100100101100;
    assign rom[1749]= 32'b11111111111111111100100011110011;
    assign rom[1750]= 32'b11111111111111111100100010111001;
    assign rom[1751]= 32'b11111111111111111100100010000000;
    assign rom[1752]= 32'b11111111111111111100100001000110;
    assign rom[1753]= 32'b11111111111111111100100000001101;
    assign rom[1754]= 32'b11111111111111111100011111010011;
    assign rom[1755]= 32'b11111111111111111100011110011010;
    assign rom[1756]= 32'b11111111111111111100011101100000;
    assign rom[1757]= 32'b11111111111111111100011100100111;
    assign rom[1758]= 32'b11111111111111111100011011101101;
    assign rom[1759]= 32'b11111111111111111100011010110011;
    assign rom[1760]= 32'b11111111111111111100011001111010;
    assign rom[1761]= 32'b11111111111111111100011001000000;
    assign rom[1762]= 32'b11111111111111111100011000000110;
    assign rom[1763]= 32'b11111111111111111100010111001101;
    assign rom[1764]= 32'b11111111111111111100010110010011;
    assign rom[1765]= 32'b11111111111111111100010101011010;
    assign rom[1766]= 32'b11111111111111111100010100100000;
    assign rom[1767]= 32'b11111111111111111100010011100111;
    assign rom[1768]= 32'b11111111111111111100010010101101;
    assign rom[1769]= 32'b11111111111111111100010001110100;
    assign rom[1770]= 32'b11111111111111111100010000111010;
    assign rom[1771]= 32'b11111111111111111100010000000001;
    assign rom[1772]= 32'b11111111111111111100001111001000;
    assign rom[1773]= 32'b11111111111111111100001110001110;
    assign rom[1774]= 32'b11111111111111111100001101010101;
    assign rom[1775]= 32'b11111111111111111100001100011100;
    assign rom[1776]= 32'b11111111111111111100001011100011;
    assign rom[1777]= 32'b11111111111111111100001010101010;
    assign rom[1778]= 32'b11111111111111111100001001110001;
    assign rom[1779]= 32'b11111111111111111100001000111000;
    assign rom[1780]= 32'b11111111111111111100000111111111;
    assign rom[1781]= 32'b11111111111111111100000111000110;
    assign rom[1782]= 32'b11111111111111111100000110001110;
    assign rom[1783]= 32'b11111111111111111100000101010101;
    assign rom[1784]= 32'b11111111111111111100000100011100;
    assign rom[1785]= 32'b11111111111111111100000011100100;
    assign rom[1786]= 32'b11111111111111111100000010101100;
    assign rom[1787]= 32'b11111111111111111100000001110100;
    assign rom[1788]= 32'b11111111111111111100000000111100;
    assign rom[1789]= 32'b11111111111111111100000000000100;
    assign rom[1790]= 32'b11111111111111111011111111001100;
    assign rom[1791]= 32'b11111111111111111011111110010100;
    assign rom[1792]= 32'b11111111111111111011111101011101;
    assign rom[1793]= 32'b11111111111111111011111100100101;
    assign rom[1794]= 32'b11111111111111111011111011101110;
    assign rom[1795]= 32'b11111111111111111011111010110111;
    assign rom[1796]= 32'b11111111111111111011111010000000;
    assign rom[1797]= 32'b11111111111111111011111001001001;
    assign rom[1798]= 32'b11111111111111111011111000010010;
    assign rom[1799]= 32'b11111111111111111011110111011100;
    assign rom[1800]= 32'b11111111111111111011110110100110;
    assign rom[1801]= 32'b11111111111111111011110101110000;
    assign rom[1802]= 32'b11111111111111111011110100111010;
    assign rom[1803]= 32'b11111111111111111011110100000100;
    assign rom[1804]= 32'b11111111111111111011110011001110;
    assign rom[1805]= 32'b11111111111111111011110010011001;
    assign rom[1806]= 32'b11111111111111111011110001100100;
    assign rom[1807]= 32'b11111111111111111011110000101111;
    assign rom[1808]= 32'b11111111111111111011101111111011;
    assign rom[1809]= 32'b11111111111111111011101111000110;
    assign rom[1810]= 32'b11111111111111111011101110010010;
    assign rom[1811]= 32'b11111111111111111011101101011110;
    assign rom[1812]= 32'b11111111111111111011101100101010;
    assign rom[1813]= 32'b11111111111111111011101011110111;
    assign rom[1814]= 32'b11111111111111111011101011000100;
    assign rom[1815]= 32'b11111111111111111011101010010001;
    assign rom[1816]= 32'b11111111111111111011101001011110;
    assign rom[1817]= 32'b11111111111111111011101000101100;
    assign rom[1818]= 32'b11111111111111111011100111111010;
    assign rom[1819]= 32'b11111111111111111011100111001000;
    assign rom[1820]= 32'b11111111111111111011100110010111;
    assign rom[1821]= 32'b11111111111111111011100101100110;
    assign rom[1822]= 32'b11111111111111111011100100110101;
    assign rom[1823]= 32'b11111111111111111011100100000100;
    assign rom[1824]= 32'b11111111111111111011100011010100;
    assign rom[1825]= 32'b11111111111111111011100010100101;
    assign rom[1826]= 32'b11111111111111111011100001110101;
    assign rom[1827]= 32'b11111111111111111011100001000110;
    assign rom[1828]= 32'b11111111111111111011100000010111;
    assign rom[1829]= 32'b11111111111111111011011111101001;
    assign rom[1830]= 32'b11111111111111111011011110111011;
    assign rom[1831]= 32'b11111111111111111011011110001101;
    assign rom[1832]= 32'b11111111111111111011011101100000;
    assign rom[1833]= 32'b11111111111111111011011100110011;
    assign rom[1834]= 32'b11111111111111111011011100000111;
    assign rom[1835]= 32'b11111111111111111011011011011011;
    assign rom[1836]= 32'b11111111111111111011011010110000;
    assign rom[1837]= 32'b11111111111111111011011010000101;
    assign rom[1838]= 32'b11111111111111111011011001011010;
    assign rom[1839]= 32'b11111111111111111011011000110000;
    assign rom[1840]= 32'b11111111111111111011011000000110;
    assign rom[1841]= 32'b11111111111111111011010111011101;
    assign rom[1842]= 32'b11111111111111111011010110110100;
    assign rom[1843]= 32'b11111111111111111011010110001100;
    assign rom[1844]= 32'b11111111111111111011010101100100;
    assign rom[1845]= 32'b11111111111111111011010100111100;
    assign rom[1846]= 32'b11111111111111111011010100010110;
    assign rom[1847]= 32'b11111111111111111011010011101111;
    assign rom[1848]= 32'b11111111111111111011010011001010;
    assign rom[1849]= 32'b11111111111111111011010010100101;
    assign rom[1850]= 32'b11111111111111111011010010000000;
    assign rom[1851]= 32'b11111111111111111011010001011100;
    assign rom[1852]= 32'b11111111111111111011010000111000;
    assign rom[1853]= 32'b11111111111111111011010000010101;
    assign rom[1854]= 32'b11111111111111111011001111110011;
    assign rom[1855]= 32'b11111111111111111011001111010001;
    assign rom[1856]= 32'b11111111111111111011001110110000;
    assign rom[1857]= 32'b11111111111111111011001110010000;
    assign rom[1858]= 32'b11111111111111111011001101110000;
    assign rom[1859]= 32'b11111111111111111011001101010001;
    assign rom[1860]= 32'b11111111111111111011001100110010;
    assign rom[1861]= 32'b11111111111111111011001100010100;
    assign rom[1862]= 32'b11111111111111111011001011110111;
    assign rom[1863]= 32'b11111111111111111011001011011010;
    assign rom[1864]= 32'b11111111111111111011001010111110;
    assign rom[1865]= 32'b11111111111111111011001010100011;
    assign rom[1866]= 32'b11111111111111111011001010001001;
    assign rom[1867]= 32'b11111111111111111011001001101111;
    assign rom[1868]= 32'b11111111111111111011001001010110;
    assign rom[1869]= 32'b11111111111111111011001000111110;
    assign rom[1870]= 32'b11111111111111111011001000100110;
    assign rom[1871]= 32'b11111111111111111011001000001111;
    assign rom[1872]= 32'b11111111111111111011000111111001;
    assign rom[1873]= 32'b11111111111111111011000111100100;
    assign rom[1874]= 32'b11111111111111111011000111010000;
    assign rom[1875]= 32'b11111111111111111011000110111100;
    assign rom[1876]= 32'b11111111111111111011000110101001;
    assign rom[1877]= 32'b11111111111111111011000110010111;
    assign rom[1878]= 32'b11111111111111111011000110000110;
    assign rom[1879]= 32'b11111111111111111011000101110110;
    assign rom[1880]= 32'b11111111111111111011000101100111;
    assign rom[1881]= 32'b11111111111111111011000101011000;
    assign rom[1882]= 32'b11111111111111111011000101001011;
    assign rom[1883]= 32'b11111111111111111011000100111110;
    assign rom[1884]= 32'b11111111111111111011000100110010;
    assign rom[1885]= 32'b11111111111111111011000100100111;
    assign rom[1886]= 32'b11111111111111111011000100011101;
    assign rom[1887]= 32'b11111111111111111011000100010100;
    assign rom[1888]= 32'b11111111111111111011000100001100;
    assign rom[1889]= 32'b11111111111111111011000100000101;
    assign rom[1890]= 32'b11111111111111111011000011111111;
    assign rom[1891]= 32'b11111111111111111011000011111010;
    assign rom[1892]= 32'b11111111111111111011000011110110;
    assign rom[1893]= 32'b11111111111111111011000011110011;
    assign rom[1894]= 32'b11111111111111111011000011110001;
    assign rom[1895]= 32'b11111111111111111011000011110000;
    assign rom[1896]= 32'b11111111111111111011000011110000;
    assign rom[1897]= 32'b11111111111111111011000011110010;
    assign rom[1898]= 32'b11111111111111111011000011110100;
    assign rom[1899]= 32'b11111111111111111011000011110111;
    assign rom[1900]= 32'b11111111111111111011000011111100;
    assign rom[1901]= 32'b11111111111111111011000100000001;
    assign rom[1902]= 32'b11111111111111111011000100001000;
    assign rom[1903]= 32'b11111111111111111011000100010000;
    assign rom[1904]= 32'b11111111111111111011000100011001;
    assign rom[1905]= 32'b11111111111111111011000100100100;
    assign rom[1906]= 32'b11111111111111111011000100101111;
    assign rom[1907]= 32'b11111111111111111011000100111100;
    assign rom[1908]= 32'b11111111111111111011000101001010;
    assign rom[1909]= 32'b11111111111111111011000101011001;
    assign rom[1910]= 32'b11111111111111111011000101101001;
    assign rom[1911]= 32'b11111111111111111011000101111011;
    assign rom[1912]= 32'b11111111111111111011000110001110;
    assign rom[1913]= 32'b11111111111111111011000110100010;
    assign rom[1914]= 32'b11111111111111111011000110111000;
    assign rom[1915]= 32'b11111111111111111011000111001110;
    assign rom[1916]= 32'b11111111111111111011000111100111;
    assign rom[1917]= 32'b11111111111111111011001000000000;
    assign rom[1918]= 32'b11111111111111111011001000011011;
    assign rom[1919]= 32'b11111111111111111011001000110111;
    assign rom[1920]= 32'b11111111111111111011001001010101;
    assign rom[1921]= 32'b11111111111111111011001001110100;
    assign rom[1922]= 32'b11111111111111111011001010010100;
    assign rom[1923]= 32'b11111111111111111011001010110110;
    assign rom[1924]= 32'b11111111111111111011001011011001;
    assign rom[1925]= 32'b11111111111111111011001011111110;
    assign rom[1926]= 32'b11111111111111111011001100100100;
    assign rom[1927]= 32'b11111111111111111011001101001100;
    assign rom[1928]= 32'b11111111111111111011001101110101;
    assign rom[1929]= 32'b11111111111111111011001110100000;
    assign rom[1930]= 32'b11111111111111111011001111001100;
    assign rom[1931]= 32'b11111111111111111011001111111010;
    assign rom[1932]= 32'b11111111111111111011010000101001;
    assign rom[1933]= 32'b11111111111111111011010001011010;
    assign rom[1934]= 32'b11111111111111111011010010001101;
    assign rom[1935]= 32'b11111111111111111011010011000001;
    assign rom[1936]= 32'b11111111111111111011010011110111;
    assign rom[1937]= 32'b11111111111111111011010100101110;
    assign rom[1938]= 32'b11111111111111111011010101100111;
    assign rom[1939]= 32'b11111111111111111011010110100001;
    assign rom[1940]= 32'b11111111111111111011010111011110;
    assign rom[1941]= 32'b11111111111111111011011000011100;
    assign rom[1942]= 32'b11111111111111111011011001011011;
    assign rom[1943]= 32'b11111111111111111011011010011101;
    assign rom[1944]= 32'b11111111111111111011011011100000;
    assign rom[1945]= 32'b11111111111111111011011100100101;
    assign rom[1946]= 32'b11111111111111111011011101101011;
    assign rom[1947]= 32'b11111111111111111011011110110011;
    assign rom[1948]= 32'b11111111111111111011011111111110;
    assign rom[1949]= 32'b11111111111111111011100001001001;
    assign rom[1950]= 32'b11111111111111111011100010010111;
    assign rom[1951]= 32'b11111111111111111011100011100111;
    assign rom[1952]= 32'b11111111111111111011100100111000;
    assign rom[1953]= 32'b11111111111111111011100110001011;
    assign rom[1954]= 32'b11111111111111111011100111100000;
    assign rom[1955]= 32'b11111111111111111011101000110111;
    assign rom[1956]= 32'b11111111111111111011101010010000;
    assign rom[1957]= 32'b11111111111111111011101011101011;
    assign rom[1958]= 32'b11111111111111111011101101001000;
    assign rom[1959]= 32'b11111111111111111011101110100110;
    assign rom[1960]= 32'b11111111111111111011110000000111;
    assign rom[1961]= 32'b11111111111111111011110001101001;
    assign rom[1962]= 32'b11111111111111111011110011001110;
    assign rom[1963]= 32'b11111111111111111011110100110100;
    assign rom[1964]= 32'b11111111111111111011110110011101;
    assign rom[1965]= 32'b11111111111111111011111000000111;
    assign rom[1966]= 32'b11111111111111111011111001110100;
    assign rom[1967]= 32'b11111111111111111011111011100010;
    assign rom[1968]= 32'b11111111111111111011111101010011;
    assign rom[1969]= 32'b11111111111111111011111111000110;
    assign rom[1970]= 32'b11111111111111111100000000111010;
    assign rom[1971]= 32'b11111111111111111100000010110001;
    assign rom[1972]= 32'b11111111111111111100000100101010;
    assign rom[1973]= 32'b11111111111111111100000110100101;
    assign rom[1974]= 32'b11111111111111111100001000100010;
    assign rom[1975]= 32'b11111111111111111100001010100010;
    assign rom[1976]= 32'b11111111111111111100001100100011;
    assign rom[1977]= 32'b11111111111111111100001110100111;
    assign rom[1978]= 32'b11111111111111111100010000101101;
    assign rom[1979]= 32'b11111111111111111100010010110101;
    assign rom[1980]= 32'b11111111111111111100010100111111;
    assign rom[1981]= 32'b11111111111111111100010111001011;
    assign rom[1982]= 32'b11111111111111111100011001011010;
    assign rom[1983]= 32'b11111111111111111100011011101011;
    assign rom[1984]= 32'b11111111111111111100011101111110;
    assign rom[1985]= 32'b11111111111111111100100000010011;
    assign rom[1986]= 32'b11111111111111111100100010101011;
    assign rom[1987]= 32'b11111111111111111100100101000101;
    assign rom[1988]= 32'b11111111111111111100100111100001;
    assign rom[1989]= 32'b11111111111111111100101001111111;
    assign rom[1990]= 32'b11111111111111111100101100100000;
    assign rom[1991]= 32'b11111111111111111100101111000011;
    assign rom[1992]= 32'b11111111111111111100110001101001;
    assign rom[1993]= 32'b11111111111111111100110100010001;
    assign rom[1994]= 32'b11111111111111111100110110111011;
    assign rom[1995]= 32'b11111111111111111100111001100111;
    assign rom[1996]= 32'b11111111111111111100111100010110;
    assign rom[1997]= 32'b11111111111111111100111111000111;
    assign rom[1998]= 32'b11111111111111111101000001111011;
    assign rom[1999]= 32'b11111111111111111101000100110001;
    assign rom[2000]= 32'b11111111111111111101000111101001;
    assign rom[2001]= 32'b11111111111111111101001010100100;
    assign rom[2002]= 32'b11111111111111111101001101100001;
    assign rom[2003]= 32'b11111111111111111101010000100001;
    assign rom[2004]= 32'b11111111111111111101010011100011;
    assign rom[2005]= 32'b11111111111111111101010110101000;
    assign rom[2006]= 32'b11111111111111111101011001101111;
    assign rom[2007]= 32'b11111111111111111101011100111000;
    assign rom[2008]= 32'b11111111111111111101100000000100;
    assign rom[2009]= 32'b11111111111111111101100011010011;
    assign rom[2010]= 32'b11111111111111111101100110100100;
    assign rom[2011]= 32'b11111111111111111101101001110111;
    assign rom[2012]= 32'b11111111111111111101101101001101;
    assign rom[2013]= 32'b11111111111111111101110000100101;
    assign rom[2014]= 32'b11111111111111111101110100000000;
    assign rom[2015]= 32'b11111111111111111101110111011110;
    assign rom[2016]= 32'b11111111111111111101111010111110;
    assign rom[2017]= 32'b11111111111111111101111110100000;
    assign rom[2018]= 32'b11111111111111111110000010000101;
    assign rom[2019]= 32'b11111111111111111110000101101101;
    assign rom[2020]= 32'b11111111111111111110001001010111;
    assign rom[2021]= 32'b11111111111111111110001101000011;
    assign rom[2022]= 32'b11111111111111111110010000110010;
    assign rom[2023]= 32'b11111111111111111110010100100100;
    assign rom[2024]= 32'b11111111111111111110011000011000;
    assign rom[2025]= 32'b11111111111111111110011100001111;
    assign rom[2026]= 32'b11111111111111111110100000001000;
    assign rom[2027]= 32'b11111111111111111110100100000100;
    assign rom[2028]= 32'b11111111111111111110101000000011;
    assign rom[2029]= 32'b11111111111111111110101100000100;
    assign rom[2030]= 32'b11111111111111111110110000000111;
    assign rom[2031]= 32'b11111111111111111110110100001110;
    assign rom[2032]= 32'b11111111111111111110111000010110;
    assign rom[2033]= 32'b11111111111111111110111100100010;
    assign rom[2034]= 32'b11111111111111111111000000110000;
    assign rom[2035]= 32'b11111111111111111111000101000000;
    assign rom[2036]= 32'b11111111111111111111001001010011;
    assign rom[2037]= 32'b11111111111111111111001101101001;
    assign rom[2038]= 32'b11111111111111111111010010000001;
    assign rom[2039]= 32'b11111111111111111111010110011100;
    assign rom[2040]= 32'b11111111111111111111011010111001;
    assign rom[2041]= 32'b11111111111111111111011111011001;
    assign rom[2042]= 32'b11111111111111111111100011111011;
    assign rom[2043]= 32'b11111111111111111111101000100001;
    assign rom[2044]= 32'b11111111111111111111101101001000;
    assign rom[2045]= 32'b11111111111111111111110001110010;
    assign rom[2046]= 32'b11111111111111111111110110011111;
    assign rom[2047]= 32'b11111111111111111111111011001111;
    assign rom[2048]= 32'b00000000000000000000000000000000;
    assign rom[2049]= 32'b00000000000000000000000100110100;
    assign rom[2050]= 32'b00000000000000000000001001101011;
    assign rom[2051]= 32'b00000000000000000000001110100101;
    assign rom[2052]= 32'b00000000000000000000010011100001;
    assign rom[2053]= 32'b00000000000000000000011000011111;
    assign rom[2054]= 32'b00000000000000000000011101100001;
    assign rom[2055]= 32'b00000000000000000000100010100100;
    assign rom[2056]= 32'b00000000000000000000100111101011;
    assign rom[2057]= 32'b00000000000000000000101100110100;
    assign rom[2058]= 32'b00000000000000000000110001111111;
    assign rom[2059]= 32'b00000000000000000000110111001101;
    assign rom[2060]= 32'b00000000000000000000111100011101;
    assign rom[2061]= 32'b00000000000000000001000001110000;
    assign rom[2062]= 32'b00000000000000000001000111000101;
    assign rom[2063]= 32'b00000000000000000001001100011101;
    assign rom[2064]= 32'b00000000000000000001010001111000;
    assign rom[2065]= 32'b00000000000000000001010111010100;
    assign rom[2066]= 32'b00000000000000000001011100110100;
    assign rom[2067]= 32'b00000000000000000001100010010101;
    assign rom[2068]= 32'b00000000000000000001100111111010;
    assign rom[2069]= 32'b00000000000000000001101101100000;
    assign rom[2070]= 32'b00000000000000000001110011001001;
    assign rom[2071]= 32'b00000000000000000001111000110101;
    assign rom[2072]= 32'b00000000000000000001111110100011;
    assign rom[2073]= 32'b00000000000000000010000100010011;
    assign rom[2074]= 32'b00000000000000000010001010000110;
    assign rom[2075]= 32'b00000000000000000010001111111011;
    assign rom[2076]= 32'b00000000000000000010010101110011;
    assign rom[2077]= 32'b00000000000000000010011011101101;
    assign rom[2078]= 32'b00000000000000000010100001101001;
    assign rom[2079]= 32'b00000000000000000010100111101000;
    assign rom[2080]= 32'b00000000000000000010101101101001;
    assign rom[2081]= 32'b00000000000000000010110011101100;
    assign rom[2082]= 32'b00000000000000000010111001110010;
    assign rom[2083]= 32'b00000000000000000010111111111001;
    assign rom[2084]= 32'b00000000000000000011000110000100;
    assign rom[2085]= 32'b00000000000000000011001100010000;
    assign rom[2086]= 32'b00000000000000000011010010011111;
    assign rom[2087]= 32'b00000000000000000011011000110000;
    assign rom[2088]= 32'b00000000000000000011011111000011;
    assign rom[2089]= 32'b00000000000000000011100101011001;
    assign rom[2090]= 32'b00000000000000000011101011110000;
    assign rom[2091]= 32'b00000000000000000011110010001010;
    assign rom[2092]= 32'b00000000000000000011111000100111;
    assign rom[2093]= 32'b00000000000000000011111111000101;
    assign rom[2094]= 32'b00000000000000000100000101100101;
    assign rom[2095]= 32'b00000000000000000100001100001000;
    assign rom[2096]= 32'b00000000000000000100010010101101;
    assign rom[2097]= 32'b00000000000000000100011001010100;
    assign rom[2098]= 32'b00000000000000000100011111111101;
    assign rom[2099]= 32'b00000000000000000100100110101000;
    assign rom[2100]= 32'b00000000000000000100101101010101;
    assign rom[2101]= 32'b00000000000000000100110100000100;
    assign rom[2102]= 32'b00000000000000000100111010110101;
    assign rom[2103]= 32'b00000000000000000101000001101001;
    assign rom[2104]= 32'b00000000000000000101001000011110;
    assign rom[2105]= 32'b00000000000000000101001111010101;
    assign rom[2106]= 32'b00000000000000000101010110001111;
    assign rom[2107]= 32'b00000000000000000101011101001010;
    assign rom[2108]= 32'b00000000000000000101100100000111;
    assign rom[2109]= 32'b00000000000000000101101011000111;
    assign rom[2110]= 32'b00000000000000000101110010001000;
    assign rom[2111]= 32'b00000000000000000101111001001011;
    assign rom[2112]= 32'b00000000000000000110000000010000;
    assign rom[2113]= 32'b00000000000000000110000111010110;
    assign rom[2114]= 32'b00000000000000000110001110011111;
    assign rom[2115]= 32'b00000000000000000110010101101001;
    assign rom[2116]= 32'b00000000000000000110011100110110;
    assign rom[2117]= 32'b00000000000000000110100100000100;
    assign rom[2118]= 32'b00000000000000000110101011010100;
    assign rom[2119]= 32'b00000000000000000110110010100101;
    assign rom[2120]= 32'b00000000000000000110111001111001;
    assign rom[2121]= 32'b00000000000000000111000001001110;
    assign rom[2122]= 32'b00000000000000000111001000100101;
    assign rom[2123]= 32'b00000000000000000111001111111101;
    assign rom[2124]= 32'b00000000000000000111010111011000;
    assign rom[2125]= 32'b00000000000000000111011110110100;
    assign rom[2126]= 32'b00000000000000000111100110010001;
    assign rom[2127]= 32'b00000000000000000111101101110000;
    assign rom[2128]= 32'b00000000000000000111110101010001;
    assign rom[2129]= 32'b00000000000000000111111100110011;
    assign rom[2130]= 32'b00000000000000001000000100010111;
    assign rom[2131]= 32'b00000000000000001000001011111101;
    assign rom[2132]= 32'b00000000000000001000010011100100;
    assign rom[2133]= 32'b00000000000000001000011011001100;
    assign rom[2134]= 32'b00000000000000001000100010110111;
    assign rom[2135]= 32'b00000000000000001000101010100010;
    assign rom[2136]= 32'b00000000000000001000110010001111;
    assign rom[2137]= 32'b00000000000000001000111001111110;
    assign rom[2138]= 32'b00000000000000001001000001101101;
    assign rom[2139]= 32'b00000000000000001001001001011111;
    assign rom[2140]= 32'b00000000000000001001010001010001;
    assign rom[2141]= 32'b00000000000000001001011001000101;
    assign rom[2142]= 32'b00000000000000001001100000111011;
    assign rom[2143]= 32'b00000000000000001001101000110010;
    assign rom[2144]= 32'b00000000000000001001110000101010;
    assign rom[2145]= 32'b00000000000000001001111000100011;
    assign rom[2146]= 32'b00000000000000001010000000011110;
    assign rom[2147]= 32'b00000000000000001010001000011010;
    assign rom[2148]= 32'b00000000000000001010010000010111;
    assign rom[2149]= 32'b00000000000000001010011000010101;
    assign rom[2150]= 32'b00000000000000001010100000010101;
    assign rom[2151]= 32'b00000000000000001010101000010101;
    assign rom[2152]= 32'b00000000000000001010110000010111;
    assign rom[2153]= 32'b00000000000000001010111000011010;
    assign rom[2154]= 32'b00000000000000001011000000011111;
    assign rom[2155]= 32'b00000000000000001011001000100100;
    assign rom[2156]= 32'b00000000000000001011010000101010;
    assign rom[2157]= 32'b00000000000000001011011000110010;
    assign rom[2158]= 32'b00000000000000001011100000111010;
    assign rom[2159]= 32'b00000000000000001011101001000100;
    assign rom[2160]= 32'b00000000000000001011110001001111;
    assign rom[2161]= 32'b00000000000000001011111001011010;
    assign rom[2162]= 32'b00000000000000001100000001100111;
    assign rom[2163]= 32'b00000000000000001100001001110101;
    assign rom[2164]= 32'b00000000000000001100010010000011;
    assign rom[2165]= 32'b00000000000000001100011010010011;
    assign rom[2166]= 32'b00000000000000001100100010100011;
    assign rom[2167]= 32'b00000000000000001100101010110101;
    assign rom[2168]= 32'b00000000000000001100110011000111;
    assign rom[2169]= 32'b00000000000000001100111011011010;
    assign rom[2170]= 32'b00000000000000001101000011101110;
    assign rom[2171]= 32'b00000000000000001101001100000011;
    assign rom[2172]= 32'b00000000000000001101010100011000;
    assign rom[2173]= 32'b00000000000000001101011100101111;
    assign rom[2174]= 32'b00000000000000001101100101000110;
    assign rom[2175]= 32'b00000000000000001101101101011110;
    assign rom[2176]= 32'b00000000000000001101110101110111;
    assign rom[2177]= 32'b00000000000000001101111110010000;
    assign rom[2178]= 32'b00000000000000001110000110101010;
    assign rom[2179]= 32'b00000000000000001110001111000101;
    assign rom[2180]= 32'b00000000000000001110010111100001;
    assign rom[2181]= 32'b00000000000000001110011111111101;
    assign rom[2182]= 32'b00000000000000001110101000011010;
    assign rom[2183]= 32'b00000000000000001110110000111000;
    assign rom[2184]= 32'b00000000000000001110111001010110;
    assign rom[2185]= 32'b00000000000000001111000001110101;
    assign rom[2186]= 32'b00000000000000001111001010010100;
    assign rom[2187]= 32'b00000000000000001111010010110100;
    assign rom[2188]= 32'b00000000000000001111011011010101;
    assign rom[2189]= 32'b00000000000000001111100011110110;
    assign rom[2190]= 32'b00000000000000001111101100010111;
    assign rom[2191]= 32'b00000000000000001111110100111001;
    assign rom[2192]= 32'b00000000000000001111111101011100;
    assign rom[2193]= 32'b00000000000000010000000101111111;
    assign rom[2194]= 32'b00000000000000010000001110100011;
    assign rom[2195]= 32'b00000000000000010000010111000111;
    assign rom[2196]= 32'b00000000000000010000011111101100;
    assign rom[2197]= 32'b00000000000000010000101000010001;
    assign rom[2198]= 32'b00000000000000010000110000110110;
    assign rom[2199]= 32'b00000000000000010000111001011100;
    assign rom[2200]= 32'b00000000000000010001000010000010;
    assign rom[2201]= 32'b00000000000000010001001010101001;
    assign rom[2202]= 32'b00000000000000010001010011010000;
    assign rom[2203]= 32'b00000000000000010001011011111000;
    assign rom[2204]= 32'b00000000000000010001100100011111;
    assign rom[2205]= 32'b00000000000000010001101101001000;
    assign rom[2206]= 32'b00000000000000010001110101110000;
    assign rom[2207]= 32'b00000000000000010001111110011001;
    assign rom[2208]= 32'b00000000000000010010000111000010;
    assign rom[2209]= 32'b00000000000000010010001111101011;
    assign rom[2210]= 32'b00000000000000010010011000010101;
    assign rom[2211]= 32'b00000000000000010010100000111111;
    assign rom[2212]= 32'b00000000000000010010101001101001;
    assign rom[2213]= 32'b00000000000000010010110010010011;
    assign rom[2214]= 32'b00000000000000010010111010111110;
    assign rom[2215]= 32'b00000000000000010011000011101001;
    assign rom[2216]= 32'b00000000000000010011001100010100;
    assign rom[2217]= 32'b00000000000000010011010100111111;
    assign rom[2218]= 32'b00000000000000010011011101101010;
    assign rom[2219]= 32'b00000000000000010011100110010110;
    assign rom[2220]= 32'b00000000000000010011101111000010;
    assign rom[2221]= 32'b00000000000000010011110111101110;
    assign rom[2222]= 32'b00000000000000010100000000011010;
    assign rom[2223]= 32'b00000000000000010100001001000110;
    assign rom[2224]= 32'b00000000000000010100010001110010;
    assign rom[2225]= 32'b00000000000000010100011010011111;
    assign rom[2226]= 32'b00000000000000010100100011001100;
    assign rom[2227]= 32'b00000000000000010100101011111000;
    assign rom[2228]= 32'b00000000000000010100110100100101;
    assign rom[2229]= 32'b00000000000000010100111101010010;
    assign rom[2230]= 32'b00000000000000010101000101111111;
    assign rom[2231]= 32'b00000000000000010101001110101100;
    assign rom[2232]= 32'b00000000000000010101010111011001;
    assign rom[2233]= 32'b00000000000000010101100000000110;
    assign rom[2234]= 32'b00000000000000010101101000110100;
    assign rom[2235]= 32'b00000000000000010101110001100001;
    assign rom[2236]= 32'b00000000000000010101111010001110;
    assign rom[2237]= 32'b00000000000000010110000010111011;
    assign rom[2238]= 32'b00000000000000010110001011101001;
    assign rom[2239]= 32'b00000000000000010110010100010110;
    assign rom[2240]= 32'b00000000000000010110011101000011;
    assign rom[2241]= 32'b00000000000000010110100101110001;
    assign rom[2242]= 32'b00000000000000010110101110011110;
    assign rom[2243]= 32'b00000000000000010110110111001011;
    assign rom[2244]= 32'b00000000000000010110111111111000;
    assign rom[2245]= 32'b00000000000000010111001000100110;
    assign rom[2246]= 32'b00000000000000010111010001010011;
    assign rom[2247]= 32'b00000000000000010111011010000000;
    assign rom[2248]= 32'b00000000000000010111100010101101;
    assign rom[2249]= 32'b00000000000000010111101011011010;
    assign rom[2250]= 32'b00000000000000010111110100000111;
    assign rom[2251]= 32'b00000000000000010111111100110100;
    assign rom[2252]= 32'b00000000000000011000000101100000;
    assign rom[2253]= 32'b00000000000000011000001110001101;
    assign rom[2254]= 32'b00000000000000011000010110111010;
    assign rom[2255]= 32'b00000000000000011000011111100110;
    assign rom[2256]= 32'b00000000000000011000101000010011;
    assign rom[2257]= 32'b00000000000000011000110000111111;
    assign rom[2258]= 32'b00000000000000011000111001101011;
    assign rom[2259]= 32'b00000000000000011001000010010111;
    assign rom[2260]= 32'b00000000000000011001001011000011;
    assign rom[2261]= 32'b00000000000000011001010011101111;
    assign rom[2262]= 32'b00000000000000011001011100011011;
    assign rom[2263]= 32'b00000000000000011001100101000110;
    assign rom[2264]= 32'b00000000000000011001101101110010;
    assign rom[2265]= 32'b00000000000000011001110110011101;
    assign rom[2266]= 32'b00000000000000011001111111001000;
    assign rom[2267]= 32'b00000000000000011010000111110011;
    assign rom[2268]= 32'b00000000000000011010010000011110;
    assign rom[2269]= 32'b00000000000000011010011001001001;
    assign rom[2270]= 32'b00000000000000011010100001110011;
    assign rom[2271]= 32'b00000000000000011010101010011110;
    assign rom[2272]= 32'b00000000000000011010110011001000;
    assign rom[2273]= 32'b00000000000000011010111011110010;
    assign rom[2274]= 32'b00000000000000011011000100011100;
    assign rom[2275]= 32'b00000000000000011011001101000101;
    assign rom[2276]= 32'b00000000000000011011010101101111;
    assign rom[2277]= 32'b00000000000000011011011110011000;
    assign rom[2278]= 32'b00000000000000011011100111000001;
    assign rom[2279]= 32'b00000000000000011011101111101010;
    assign rom[2280]= 32'b00000000000000011011111000010011;
    assign rom[2281]= 32'b00000000000000011100000000111100;
    assign rom[2282]= 32'b00000000000000011100001001100100;
    assign rom[2283]= 32'b00000000000000011100010010001100;
    assign rom[2284]= 32'b00000000000000011100011010110100;
    assign rom[2285]= 32'b00000000000000011100100011011100;
    assign rom[2286]= 32'b00000000000000011100101100000100;
    assign rom[2287]= 32'b00000000000000011100110100101011;
    assign rom[2288]= 32'b00000000000000011100111101010010;
    assign rom[2289]= 32'b00000000000000011101000101111001;
    assign rom[2290]= 32'b00000000000000011101001110100000;
    assign rom[2291]= 32'b00000000000000011101010111000110;
    assign rom[2292]= 32'b00000000000000011101011111101101;
    assign rom[2293]= 32'b00000000000000011101101000010011;
    assign rom[2294]= 32'b00000000000000011101110000111000;
    assign rom[2295]= 32'b00000000000000011101111001011110;
    assign rom[2296]= 32'b00000000000000011110000010000100;
    assign rom[2297]= 32'b00000000000000011110001010101001;
    assign rom[2298]= 32'b00000000000000011110010011001110;
    assign rom[2299]= 32'b00000000000000011110011011110010;
    assign rom[2300]= 32'b00000000000000011110100100010111;
    assign rom[2301]= 32'b00000000000000011110101100111011;
    assign rom[2302]= 32'b00000000000000011110110101011111;
    assign rom[2303]= 32'b00000000000000011110111110000011;
    assign rom[2304]= 32'b00000000000000011111000110100111;
    assign rom[2305]= 32'b00000000000000011111001111001010;
    assign rom[2306]= 32'b00000000000000011111010111101101;
    assign rom[2307]= 32'b00000000000000011111100000010000;
    assign rom[2308]= 32'b00000000000000011111101000110011;
    assign rom[2309]= 32'b00000000000000011111110001010101;
    assign rom[2310]= 32'b00000000000000011111111001111000;
    assign rom[2311]= 32'b00000000000000100000000010011010;
    assign rom[2312]= 32'b00000000000000100000001010111011;
    assign rom[2313]= 32'b00000000000000100000010011011101;
    assign rom[2314]= 32'b00000000000000100000011011111110;
    assign rom[2315]= 32'b00000000000000100000100100011111;
    assign rom[2316]= 32'b00000000000000100000101101000000;
    assign rom[2317]= 32'b00000000000000100000110101100000;
    assign rom[2318]= 32'b00000000000000100000111110000001;
    assign rom[2319]= 32'b00000000000000100001000110100001;
    assign rom[2320]= 32'b00000000000000100001001111000001;
    assign rom[2321]= 32'b00000000000000100001010111100000;
    assign rom[2322]= 32'b00000000000000100001100000000000;
    assign rom[2323]= 32'b00000000000000100001101000011111;
    assign rom[2324]= 32'b00000000000000100001110000111110;
    assign rom[2325]= 32'b00000000000000100001111001011100;
    assign rom[2326]= 32'b00000000000000100010000001111011;
    assign rom[2327]= 32'b00000000000000100010001010011001;
    assign rom[2328]= 32'b00000000000000100010010010110111;
    assign rom[2329]= 32'b00000000000000100010011011010101;
    assign rom[2330]= 32'b00000000000000100010100011110010;
    assign rom[2331]= 32'b00000000000000100010101100010000;
    assign rom[2332]= 32'b00000000000000100010110100101101;
    assign rom[2333]= 32'b00000000000000100010111101001001;
    assign rom[2334]= 32'b00000000000000100011000101100110;
    assign rom[2335]= 32'b00000000000000100011001110000010;
    assign rom[2336]= 32'b00000000000000100011010110011110;
    assign rom[2337]= 32'b00000000000000100011011110111010;
    assign rom[2338]= 32'b00000000000000100011100111010110;
    assign rom[2339]= 32'b00000000000000100011101111110001;
    assign rom[2340]= 32'b00000000000000100011111000001101;
    assign rom[2341]= 32'b00000000000000100100000000101000;
    assign rom[2342]= 32'b00000000000000100100001001000010;
    assign rom[2343]= 32'b00000000000000100100010001011101;
    assign rom[2344]= 32'b00000000000000100100011001110111;
    assign rom[2345]= 32'b00000000000000100100100010010001;
    assign rom[2346]= 32'b00000000000000100100101010101011;
    assign rom[2347]= 32'b00000000000000100100110011000101;
    assign rom[2348]= 32'b00000000000000100100111011011110;
    assign rom[2349]= 32'b00000000000000100101000011110111;
    assign rom[2350]= 32'b00000000000000100101001100010000;
    assign rom[2351]= 32'b00000000000000100101010100101001;
    assign rom[2352]= 32'b00000000000000100101011101000001;
    assign rom[2353]= 32'b00000000000000100101100101011010;
    assign rom[2354]= 32'b00000000000000100101101101110010;
    assign rom[2355]= 32'b00000000000000100101110110001010;
    assign rom[2356]= 32'b00000000000000100101111110100001;
    assign rom[2357]= 32'b00000000000000100110000110111001;
    assign rom[2358]= 32'b00000000000000100110001111010000;
    assign rom[2359]= 32'b00000000000000100110010111100111;
    assign rom[2360]= 32'b00000000000000100110011111111110;
    assign rom[2361]= 32'b00000000000000100110101000010100;
    assign rom[2362]= 32'b00000000000000100110110000101011;
    assign rom[2363]= 32'b00000000000000100110111001000001;
    assign rom[2364]= 32'b00000000000000100111000001010111;
    assign rom[2365]= 32'b00000000000000100111001001101101;
    assign rom[2366]= 32'b00000000000000100111010010000010;
    assign rom[2367]= 32'b00000000000000100111011010011000;
    assign rom[2368]= 32'b00000000000000100111100010101101;
    assign rom[2369]= 32'b00000000000000100111101011000010;
    assign rom[2370]= 32'b00000000000000100111110011010110;
    assign rom[2371]= 32'b00000000000000100111111011101011;
    assign rom[2372]= 32'b00000000000000101000000011111111;
    assign rom[2373]= 32'b00000000000000101000001100010011;
    assign rom[2374]= 32'b00000000000000101000010100100111;
    assign rom[2375]= 32'b00000000000000101000011100111011;
    assign rom[2376]= 32'b00000000000000101000100101001111;
    assign rom[2377]= 32'b00000000000000101000101101100010;
    assign rom[2378]= 32'b00000000000000101000110101110101;
    assign rom[2379]= 32'b00000000000000101000111110001000;
    assign rom[2380]= 32'b00000000000000101001000110011011;
    assign rom[2381]= 32'b00000000000000101001001110101110;
    assign rom[2382]= 32'b00000000000000101001010111000000;
    assign rom[2383]= 32'b00000000000000101001011111010011;
    assign rom[2384]= 32'b00000000000000101001100111100101;
    assign rom[2385]= 32'b00000000000000101001101111110111;
    assign rom[2386]= 32'b00000000000000101001111000001000;
    assign rom[2387]= 32'b00000000000000101010000000011010;
    assign rom[2388]= 32'b00000000000000101010001000101011;
    assign rom[2389]= 32'b00000000000000101010010000111101;
    assign rom[2390]= 32'b00000000000000101010011001001110;
    assign rom[2391]= 32'b00000000000000101010100001011111;
    assign rom[2392]= 32'b00000000000000101010101001101111;
    assign rom[2393]= 32'b00000000000000101010110010000000;
    assign rom[2394]= 32'b00000000000000101010111010010000;
    assign rom[2395]= 32'b00000000000000101011000010100000;
    assign rom[2396]= 32'b00000000000000101011001010110000;
    assign rom[2397]= 32'b00000000000000101011010011000000;
    assign rom[2398]= 32'b00000000000000101011011011010000;
    assign rom[2399]= 32'b00000000000000101011100011011111;
    assign rom[2400]= 32'b00000000000000101011101011101111;
    assign rom[2401]= 32'b00000000000000101011110011111110;
    assign rom[2402]= 32'b00000000000000101011111100001101;
    assign rom[2403]= 32'b00000000000000101100000100011100;
    assign rom[2404]= 32'b00000000000000101100001100101011;
    assign rom[2405]= 32'b00000000000000101100010100111001;
    assign rom[2406]= 32'b00000000000000101100011101001000;
    assign rom[2407]= 32'b00000000000000101100100101010110;
    assign rom[2408]= 32'b00000000000000101100101101100100;
    assign rom[2409]= 32'b00000000000000101100110101110010;
    assign rom[2410]= 32'b00000000000000101100111110000000;
    assign rom[2411]= 32'b00000000000000101101000110001110;
    assign rom[2412]= 32'b00000000000000101101001110011011;
    assign rom[2413]= 32'b00000000000000101101010110101001;
    assign rom[2414]= 32'b00000000000000101101011110110110;
    assign rom[2415]= 32'b00000000000000101101100111000011;
    assign rom[2416]= 32'b00000000000000101101101111010000;
    assign rom[2417]= 32'b00000000000000101101110111011101;
    assign rom[2418]= 32'b00000000000000101101111111101001;
    assign rom[2419]= 32'b00000000000000101110000111110110;
    assign rom[2420]= 32'b00000000000000101110010000000010;
    assign rom[2421]= 32'b00000000000000101110011000001111;
    assign rom[2422]= 32'b00000000000000101110100000011011;
    assign rom[2423]= 32'b00000000000000101110101000100111;
    assign rom[2424]= 32'b00000000000000101110110000110011;
    assign rom[2425]= 32'b00000000000000101110111000111110;
    assign rom[2426]= 32'b00000000000000101111000001001010;
    assign rom[2427]= 32'b00000000000000101111001001010101;
    assign rom[2428]= 32'b00000000000000101111010001100001;
    assign rom[2429]= 32'b00000000000000101111011001101100;
    assign rom[2430]= 32'b00000000000000101111100001110111;
    assign rom[2431]= 32'b00000000000000101111101010000010;
    assign rom[2432]= 32'b00000000000000101111110010001101;
    assign rom[2433]= 32'b00000000000000101111111010011000;
    assign rom[2434]= 32'b00000000000000110000000010100010;
    assign rom[2435]= 32'b00000000000000110000001010101101;
    assign rom[2436]= 32'b00000000000000110000010010110111;
    assign rom[2437]= 32'b00000000000000110000011011000010;
    assign rom[2438]= 32'b00000000000000110000100011001100;
    assign rom[2439]= 32'b00000000000000110000101011010110;
    assign rom[2440]= 32'b00000000000000110000110011100000;
    assign rom[2441]= 32'b00000000000000110000111011101010;
    assign rom[2442]= 32'b00000000000000110001000011110011;
    assign rom[2443]= 32'b00000000000000110001001011111101;
    assign rom[2444]= 32'b00000000000000110001010100000110;
    assign rom[2445]= 32'b00000000000000110001011100010000;
    assign rom[2446]= 32'b00000000000000110001100100011001;
    assign rom[2447]= 32'b00000000000000110001101100100010;
    assign rom[2448]= 32'b00000000000000110001110100101011;
    assign rom[2449]= 32'b00000000000000110001111100110100;
    assign rom[2450]= 32'b00000000000000110010000100111101;
    assign rom[2451]= 32'b00000000000000110010001101000110;
    assign rom[2452]= 32'b00000000000000110010010101001110;
    assign rom[2453]= 32'b00000000000000110010011101010111;
    assign rom[2454]= 32'b00000000000000110010100101011111;
    assign rom[2455]= 32'b00000000000000110010101101101000;
    assign rom[2456]= 32'b00000000000000110010110101110000;
    assign rom[2457]= 32'b00000000000000110010111101111000;
    assign rom[2458]= 32'b00000000000000110011000110000000;
    assign rom[2459]= 32'b00000000000000110011001110001000;
    assign rom[2460]= 32'b00000000000000110011010110010000;
    assign rom[2461]= 32'b00000000000000110011011110011000;
    assign rom[2462]= 32'b00000000000000110011100110100000;
    assign rom[2463]= 32'b00000000000000110011101110100111;
    assign rom[2464]= 32'b00000000000000110011110110101111;
    assign rom[2465]= 32'b00000000000000110011111110110110;
    assign rom[2466]= 32'b00000000000000110100000110111110;
    assign rom[2467]= 32'b00000000000000110100001111000101;
    assign rom[2468]= 32'b00000000000000110100010111001100;
    assign rom[2469]= 32'b00000000000000110100011111010011;
    assign rom[2470]= 32'b00000000000000110100100111011010;
    assign rom[2471]= 32'b00000000000000110100101111100001;
    assign rom[2472]= 32'b00000000000000110100110111101000;
    assign rom[2473]= 32'b00000000000000110100111111101111;
    assign rom[2474]= 32'b00000000000000110101000111110101;
    assign rom[2475]= 32'b00000000000000110101001111111100;
    assign rom[2476]= 32'b00000000000000110101011000000010;
    assign rom[2477]= 32'b00000000000000110101100000001001;
    assign rom[2478]= 32'b00000000000000110101101000001111;
    assign rom[2479]= 32'b00000000000000110101110000010110;
    assign rom[2480]= 32'b00000000000000110101111000011100;
    assign rom[2481]= 32'b00000000000000110110000000100010;
    assign rom[2482]= 32'b00000000000000110110001000101000;
    assign rom[2483]= 32'b00000000000000110110010000101110;
    assign rom[2484]= 32'b00000000000000110110011000110100;
    assign rom[2485]= 32'b00000000000000110110100000111010;
    assign rom[2486]= 32'b00000000000000110110101001000000;
    assign rom[2487]= 32'b00000000000000110110110001000101;
    assign rom[2488]= 32'b00000000000000110110111001001011;
    assign rom[2489]= 32'b00000000000000110111000001010000;
    assign rom[2490]= 32'b00000000000000110111001001010110;
    assign rom[2491]= 32'b00000000000000110111010001011011;
    assign rom[2492]= 32'b00000000000000110111011001100001;
    assign rom[2493]= 32'b00000000000000110111100001100110;
    assign rom[2494]= 32'b00000000000000110111101001101011;
    assign rom[2495]= 32'b00000000000000110111110001110001;
    assign rom[2496]= 32'b00000000000000110111111001110110;
    assign rom[2497]= 32'b00000000000000111000000001111011;
    assign rom[2498]= 32'b00000000000000111000001010000000;
    assign rom[2499]= 32'b00000000000000111000010010000101;
    assign rom[2500]= 32'b00000000000000111000011010001010;
    assign rom[2501]= 32'b00000000000000111000100010001110;
    assign rom[2502]= 32'b00000000000000111000101010010011;
    assign rom[2503]= 32'b00000000000000111000110010011000;
    assign rom[2504]= 32'b00000000000000111000111010011100;
    assign rom[2505]= 32'b00000000000000111001000010100001;
    assign rom[2506]= 32'b00000000000000111001001010100110;
    assign rom[2507]= 32'b00000000000000111001010010101010;
    assign rom[2508]= 32'b00000000000000111001011010101110;
    assign rom[2509]= 32'b00000000000000111001100010110011;
    assign rom[2510]= 32'b00000000000000111001101010110111;
    assign rom[2511]= 32'b00000000000000111001110010111011;
    assign rom[2512]= 32'b00000000000000111001111011000000;
    assign rom[2513]= 32'b00000000000000111010000011000100;
    assign rom[2514]= 32'b00000000000000111010001011001000;
    assign rom[2515]= 32'b00000000000000111010010011001100;
    assign rom[2516]= 32'b00000000000000111010011011010000;
    assign rom[2517]= 32'b00000000000000111010100011010100;
    assign rom[2518]= 32'b00000000000000111010101011011000;
    assign rom[2519]= 32'b00000000000000111010110011011100;
    assign rom[2520]= 32'b00000000000000111010111011011111;
    assign rom[2521]= 32'b00000000000000111011000011100011;
    assign rom[2522]= 32'b00000000000000111011001011100111;
    assign rom[2523]= 32'b00000000000000111011010011101010;
    assign rom[2524]= 32'b00000000000000111011011011101110;
    assign rom[2525]= 32'b00000000000000111011100011110010;
    assign rom[2526]= 32'b00000000000000111011101011110101;
    assign rom[2527]= 32'b00000000000000111011110011111001;
    assign rom[2528]= 32'b00000000000000111011111011111100;
    assign rom[2529]= 32'b00000000000000111100000100000000;
    assign rom[2530]= 32'b00000000000000111100001100000011;
    assign rom[2531]= 32'b00000000000000111100010100000110;
    assign rom[2532]= 32'b00000000000000111100011100001001;
    assign rom[2533]= 32'b00000000000000111100100100001101;
    assign rom[2534]= 32'b00000000000000111100101100010000;
    assign rom[2535]= 32'b00000000000000111100110100010011;
    assign rom[2536]= 32'b00000000000000111100111100010110;
    assign rom[2537]= 32'b00000000000000111101000100011001;
    assign rom[2538]= 32'b00000000000000111101001100011100;
    assign rom[2539]= 32'b00000000000000111101010100011111;
    assign rom[2540]= 32'b00000000000000111101011100100010;
    assign rom[2541]= 32'b00000000000000111101100100100101;
    assign rom[2542]= 32'b00000000000000111101101100101000;
    assign rom[2543]= 32'b00000000000000111101110100101011;
    assign rom[2544]= 32'b00000000000000111101111100101110;
    assign rom[2545]= 32'b00000000000000111110000100110000;
    assign rom[2546]= 32'b00000000000000111110001100110011;
    assign rom[2547]= 32'b00000000000000111110010100110110;
    assign rom[2548]= 32'b00000000000000111110011100111000;
    assign rom[2549]= 32'b00000000000000111110100100111011;
    assign rom[2550]= 32'b00000000000000111110101100111110;
    assign rom[2551]= 32'b00000000000000111110110101000000;
    assign rom[2552]= 32'b00000000000000111110111101000011;
    assign rom[2553]= 32'b00000000000000111111000101000101;
    assign rom[2554]= 32'b00000000000000111111001101001000;
    assign rom[2555]= 32'b00000000000000111111010101001010;
    assign rom[2556]= 32'b00000000000000111111011101001101;
    assign rom[2557]= 32'b00000000000000111111100101001111;
    assign rom[2558]= 32'b00000000000000111111101101010001;
    assign rom[2559]= 32'b00000000000000111111110101010100;
    assign rom[2560]= 32'b00000000000000111111111101010110;
    assign rom[2561]= 32'b00000000000001000000000101011000;
    assign rom[2562]= 32'b00000000000001000000001101011010;
    assign rom[2563]= 32'b00000000000001000000010101011101;
    assign rom[2564]= 32'b00000000000001000000011101011111;
    assign rom[2565]= 32'b00000000000001000000100101100001;
    assign rom[2566]= 32'b00000000000001000000101101100011;
    assign rom[2567]= 32'b00000000000001000000110101100101;
    assign rom[2568]= 32'b00000000000001000000111101100111;
    assign rom[2569]= 32'b00000000000001000001000101101001;
    assign rom[2570]= 32'b00000000000001000001001101101011;
    assign rom[2571]= 32'b00000000000001000001010101101101;
    assign rom[2572]= 32'b00000000000001000001011101101111;
    assign rom[2573]= 32'b00000000000001000001100101110001;
    assign rom[2574]= 32'b00000000000001000001101101110011;
    assign rom[2575]= 32'b00000000000001000001110101110101;
    assign rom[2576]= 32'b00000000000001000001111101110111;
    assign rom[2577]= 32'b00000000000001000010000101111001;
    assign rom[2578]= 32'b00000000000001000010001101111010;
    assign rom[2579]= 32'b00000000000001000010010101111100;
    assign rom[2580]= 32'b00000000000001000010011101111110;
    assign rom[2581]= 32'b00000000000001000010100110000000;
    assign rom[2582]= 32'b00000000000001000010101110000001;
    assign rom[2583]= 32'b00000000000001000010110110000011;
    assign rom[2584]= 32'b00000000000001000010111110000101;
    assign rom[2585]= 32'b00000000000001000011000110000110;
    assign rom[2586]= 32'b00000000000001000011001110001000;
    assign rom[2587]= 32'b00000000000001000011010110001010;
    assign rom[2588]= 32'b00000000000001000011011110001011;
    assign rom[2589]= 32'b00000000000001000011100110001101;
    assign rom[2590]= 32'b00000000000001000011101110001110;
    assign rom[2591]= 32'b00000000000001000011110110010000;
    assign rom[2592]= 32'b00000000000001000011111110010001;
    assign rom[2593]= 32'b00000000000001000100000110010011;
    assign rom[2594]= 32'b00000000000001000100001110010100;
    assign rom[2595]= 32'b00000000000001000100010110010110;
    assign rom[2596]= 32'b00000000000001000100011110010111;
    assign rom[2597]= 32'b00000000000001000100100110011001;
    assign rom[2598]= 32'b00000000000001000100101110011010;
    assign rom[2599]= 32'b00000000000001000100110110011011;
    assign rom[2600]= 32'b00000000000001000100111110011101;
    assign rom[2601]= 32'b00000000000001000101000110011110;
    assign rom[2602]= 32'b00000000000001000101001110011111;
    assign rom[2603]= 32'b00000000000001000101010110100001;
    assign rom[2604]= 32'b00000000000001000101011110100010;
    assign rom[2605]= 32'b00000000000001000101100110100011;
    assign rom[2606]= 32'b00000000000001000101101110100100;
    assign rom[2607]= 32'b00000000000001000101110110100110;
    assign rom[2608]= 32'b00000000000001000101111110100111;
    assign rom[2609]= 32'b00000000000001000110000110101000;
    assign rom[2610]= 32'b00000000000001000110001110101001;
    assign rom[2611]= 32'b00000000000001000110010110101010;
    assign rom[2612]= 32'b00000000000001000110011110101100;
    assign rom[2613]= 32'b00000000000001000110100110101101;
    assign rom[2614]= 32'b00000000000001000110101110101110;
    assign rom[2615]= 32'b00000000000001000110110110101111;
    assign rom[2616]= 32'b00000000000001000110111110110000;
    assign rom[2617]= 32'b00000000000001000111000110110001;
    assign rom[2618]= 32'b00000000000001000111001110110010;
    assign rom[2619]= 32'b00000000000001000111010110110011;
    assign rom[2620]= 32'b00000000000001000111011110110100;
    assign rom[2621]= 32'b00000000000001000111100110110101;
    assign rom[2622]= 32'b00000000000001000111101110110110;
    assign rom[2623]= 32'b00000000000001000111110110110111;
    assign rom[2624]= 32'b00000000000001000111111110111000;
    assign rom[2625]= 32'b00000000000001001000000110111001;
    assign rom[2626]= 32'b00000000000001001000001110111010;
    assign rom[2627]= 32'b00000000000001001000010110111011;
    assign rom[2628]= 32'b00000000000001001000011110111100;
    assign rom[2629]= 32'b00000000000001001000100110111101;
    assign rom[2630]= 32'b00000000000001001000101110111110;
    assign rom[2631]= 32'b00000000000001001000110110111111;
    assign rom[2632]= 32'b00000000000001001000111111000000;
    assign rom[2633]= 32'b00000000000001001001000111000001;
    assign rom[2634]= 32'b00000000000001001001001111000001;
    assign rom[2635]= 32'b00000000000001001001010111000010;
    assign rom[2636]= 32'b00000000000001001001011111000011;
    assign rom[2637]= 32'b00000000000001001001100111000100;
    assign rom[2638]= 32'b00000000000001001001101111000101;
    assign rom[2639]= 32'b00000000000001001001110111000110;
    assign rom[2640]= 32'b00000000000001001001111111000110;
    assign rom[2641]= 32'b00000000000001001010000111000111;
    assign rom[2642]= 32'b00000000000001001010001111001000;
    assign rom[2643]= 32'b00000000000001001010010111001001;
    assign rom[2644]= 32'b00000000000001001010011111001001;
    assign rom[2645]= 32'b00000000000001001010100111001010;
    assign rom[2646]= 32'b00000000000001001010101111001011;
    assign rom[2647]= 32'b00000000000001001010110111001100;
    assign rom[2648]= 32'b00000000000001001010111111001100;
    assign rom[2649]= 32'b00000000000001001011000111001101;
    assign rom[2650]= 32'b00000000000001001011001111001110;
    assign rom[2651]= 32'b00000000000001001011010111001110;
    assign rom[2652]= 32'b00000000000001001011011111001111;
    assign rom[2653]= 32'b00000000000001001011100111010000;
    assign rom[2654]= 32'b00000000000001001011101111010000;
    assign rom[2655]= 32'b00000000000001001011110111010001;
    assign rom[2656]= 32'b00000000000001001011111111010010;
    assign rom[2657]= 32'b00000000000001001100000111010010;
    assign rom[2658]= 32'b00000000000001001100001111010011;
    assign rom[2659]= 32'b00000000000001001100010111010100;
    assign rom[2660]= 32'b00000000000001001100011111010100;
    assign rom[2661]= 32'b00000000000001001100100111010101;
    assign rom[2662]= 32'b00000000000001001100101111010101;
    assign rom[2663]= 32'b00000000000001001100110111010110;
    assign rom[2664]= 32'b00000000000001001100111111010111;
    assign rom[2665]= 32'b00000000000001001101000111010111;
    assign rom[2666]= 32'b00000000000001001101001111011000;
    assign rom[2667]= 32'b00000000000001001101010111011000;
    assign rom[2668]= 32'b00000000000001001101011111011001;
    assign rom[2669]= 32'b00000000000001001101100111011001;
    assign rom[2670]= 32'b00000000000001001101101111011010;
    assign rom[2671]= 32'b00000000000001001101110111011010;
    assign rom[2672]= 32'b00000000000001001101111111011011;
    assign rom[2673]= 32'b00000000000001001110000111011011;
    assign rom[2674]= 32'b00000000000001001110001111011100;
    assign rom[2675]= 32'b00000000000001001110010111011100;
    assign rom[2676]= 32'b00000000000001001110011111011101;
    assign rom[2677]= 32'b00000000000001001110100111011101;
    assign rom[2678]= 32'b00000000000001001110101111011110;
    assign rom[2679]= 32'b00000000000001001110110111011110;
    assign rom[2680]= 32'b00000000000001001110111111011111;
    assign rom[2681]= 32'b00000000000001001111000111011111;
    assign rom[2682]= 32'b00000000000001001111001111100000;
    assign rom[2683]= 32'b00000000000001001111010111100000;
    assign rom[2684]= 32'b00000000000001001111011111100000;
    assign rom[2685]= 32'b00000000000001001111100111100001;
    assign rom[2686]= 32'b00000000000001001111101111100001;
    assign rom[2687]= 32'b00000000000001001111110111100010;
    assign rom[2688]= 32'b00000000000001001111111111100010;
    assign rom[2689]= 32'b00000000000001010000000111100011;
    assign rom[2690]= 32'b00000000000001010000001111100011;
    assign rom[2691]= 32'b00000000000001010000010111100011;
    assign rom[2692]= 32'b00000000000001010000011111100100;
    assign rom[2693]= 32'b00000000000001010000100111100100;
    assign rom[2694]= 32'b00000000000001010000101111100101;
    assign rom[2695]= 32'b00000000000001010000110111100101;
    assign rom[2696]= 32'b00000000000001010000111111100101;
    assign rom[2697]= 32'b00000000000001010001000111100110;
    assign rom[2698]= 32'b00000000000001010001001111100110;
    assign rom[2699]= 32'b00000000000001010001010111100110;
    assign rom[2700]= 32'b00000000000001010001011111100111;
    assign rom[2701]= 32'b00000000000001010001100111100111;
    assign rom[2702]= 32'b00000000000001010001101111100111;
    assign rom[2703]= 32'b00000000000001010001110111101000;
    assign rom[2704]= 32'b00000000000001010001111111101000;
    assign rom[2705]= 32'b00000000000001010010000111101000;
    assign rom[2706]= 32'b00000000000001010010001111101001;
    assign rom[2707]= 32'b00000000000001010010010111101001;
    assign rom[2708]= 32'b00000000000001010010011111101001;
    assign rom[2709]= 32'b00000000000001010010100111101010;
    assign rom[2710]= 32'b00000000000001010010101111101010;
    assign rom[2711]= 32'b00000000000001010010110111101010;
    assign rom[2712]= 32'b00000000000001010010111111101011;
    assign rom[2713]= 32'b00000000000001010011000111101011;
    assign rom[2714]= 32'b00000000000001010011001111101011;
    assign rom[2715]= 32'b00000000000001010011010111101011;
    assign rom[2716]= 32'b00000000000001010011011111101100;
    assign rom[2717]= 32'b00000000000001010011100111101100;
    assign rom[2718]= 32'b00000000000001010011101111101100;
    assign rom[2719]= 32'b00000000000001010011110111101100;
    assign rom[2720]= 32'b00000000000001010011111111101101;
    assign rom[2721]= 32'b00000000000001010100000111101101;
    assign rom[2722]= 32'b00000000000001010100001111101101;
    assign rom[2723]= 32'b00000000000001010100010111101110;
    assign rom[2724]= 32'b00000000000001010100011111101110;
    assign rom[2725]= 32'b00000000000001010100100111101110;
    assign rom[2726]= 32'b00000000000001010100101111101110;
    assign rom[2727]= 32'b00000000000001010100110111101111;
    assign rom[2728]= 32'b00000000000001010100111111101111;
    assign rom[2729]= 32'b00000000000001010101000111101111;
    assign rom[2730]= 32'b00000000000001010101001111101111;
    assign rom[2731]= 32'b00000000000001010101010111101111;
    assign rom[2732]= 32'b00000000000001010101011111110000;
    assign rom[2733]= 32'b00000000000001010101100111110000;
    assign rom[2734]= 32'b00000000000001010101101111110000;
    assign rom[2735]= 32'b00000000000001010101110111110000;
    assign rom[2736]= 32'b00000000000001010101111111110001;
    assign rom[2737]= 32'b00000000000001010110000111110001;
    assign rom[2738]= 32'b00000000000001010110001111110001;
    assign rom[2739]= 32'b00000000000001010110010111110001;
    assign rom[2740]= 32'b00000000000001010110011111110001;
    assign rom[2741]= 32'b00000000000001010110100111110010;
    assign rom[2742]= 32'b00000000000001010110101111110010;
    assign rom[2743]= 32'b00000000000001010110110111110010;
    assign rom[2744]= 32'b00000000000001010110111111110010;
    assign rom[2745]= 32'b00000000000001010111000111110010;
    assign rom[2746]= 32'b00000000000001010111001111110011;
    assign rom[2747]= 32'b00000000000001010111010111110011;
    assign rom[2748]= 32'b00000000000001010111011111110011;
    assign rom[2749]= 32'b00000000000001010111100111110011;
    assign rom[2750]= 32'b00000000000001010111101111110011;
    assign rom[2751]= 32'b00000000000001010111110111110011;
    assign rom[2752]= 32'b00000000000001010111111111110100;
    assign rom[2753]= 32'b00000000000001011000000111110100;
    assign rom[2754]= 32'b00000000000001011000001111110100;
    assign rom[2755]= 32'b00000000000001011000010111110100;
    assign rom[2756]= 32'b00000000000001011000011111110100;
    assign rom[2757]= 32'b00000000000001011000100111110100;
    assign rom[2758]= 32'b00000000000001011000101111110101;
    assign rom[2759]= 32'b00000000000001011000110111110101;
    assign rom[2760]= 32'b00000000000001011000111111110101;
    assign rom[2761]= 32'b00000000000001011001000111110101;
    assign rom[2762]= 32'b00000000000001011001001111110101;
    assign rom[2763]= 32'b00000000000001011001010111110101;
    assign rom[2764]= 32'b00000000000001011001011111110101;
    assign rom[2765]= 32'b00000000000001011001100111110110;
    assign rom[2766]= 32'b00000000000001011001101111110110;
    assign rom[2767]= 32'b00000000000001011001110111110110;
    assign rom[2768]= 32'b00000000000001011001111111110110;
    assign rom[2769]= 32'b00000000000001011010000111110110;
    assign rom[2770]= 32'b00000000000001011010001111110110;
    assign rom[2771]= 32'b00000000000001011010010111110110;
    assign rom[2772]= 32'b00000000000001011010011111110111;
    assign rom[2773]= 32'b00000000000001011010100111110111;
    assign rom[2774]= 32'b00000000000001011010101111110111;
    assign rom[2775]= 32'b00000000000001011010110111110111;
    assign rom[2776]= 32'b00000000000001011010111111110111;
    assign rom[2777]= 32'b00000000000001011011000111110111;
    assign rom[2778]= 32'b00000000000001011011001111110111;
    assign rom[2779]= 32'b00000000000001011011010111110111;
    assign rom[2780]= 32'b00000000000001011011011111110111;
    assign rom[2781]= 32'b00000000000001011011100111111000;
    assign rom[2782]= 32'b00000000000001011011101111111000;
    assign rom[2783]= 32'b00000000000001011011110111111000;
    assign rom[2784]= 32'b00000000000001011011111111111000;
    assign rom[2785]= 32'b00000000000001011100000111111000;
    assign rom[2786]= 32'b00000000000001011100001111111000;
    assign rom[2787]= 32'b00000000000001011100010111111000;
    assign rom[2788]= 32'b00000000000001011100011111111000;
    assign rom[2789]= 32'b00000000000001011100100111111000;
    assign rom[2790]= 32'b00000000000001011100101111111001;
    assign rom[2791]= 32'b00000000000001011100110111111001;
    assign rom[2792]= 32'b00000000000001011100111111111001;
    assign rom[2793]= 32'b00000000000001011101000111111001;
    assign rom[2794]= 32'b00000000000001011101001111111001;
    assign rom[2795]= 32'b00000000000001011101010111111001;
    assign rom[2796]= 32'b00000000000001011101011111111001;
    assign rom[2797]= 32'b00000000000001011101100111111001;
    assign rom[2798]= 32'b00000000000001011101101111111001;
    assign rom[2799]= 32'b00000000000001011101110111111001;
    assign rom[2800]= 32'b00000000000001011101111111111001;
    assign rom[2801]= 32'b00000000000001011110000111111010;
    assign rom[2802]= 32'b00000000000001011110001111111010;
    assign rom[2803]= 32'b00000000000001011110010111111010;
    assign rom[2804]= 32'b00000000000001011110011111111010;
    assign rom[2805]= 32'b00000000000001011110100111111010;
    assign rom[2806]= 32'b00000000000001011110101111111010;
    assign rom[2807]= 32'b00000000000001011110110111111010;
    assign rom[2808]= 32'b00000000000001011110111111111010;
    assign rom[2809]= 32'b00000000000001011111000111111010;
    assign rom[2810]= 32'b00000000000001011111001111111010;
    assign rom[2811]= 32'b00000000000001011111010111111010;
    assign rom[2812]= 32'b00000000000001011111011111111010;
    assign rom[2813]= 32'b00000000000001011111100111111010;
    assign rom[2814]= 32'b00000000000001011111101111111011;
    assign rom[2815]= 32'b00000000000001011111110111111011;
    assign rom[2816]= 32'b00000000000001011111111111111011;
    assign rom[2817]= 32'b00000000000001100000000111111011;
    assign rom[2818]= 32'b00000000000001100000001111111011;
    assign rom[2819]= 32'b00000000000001100000010111111011;
    assign rom[2820]= 32'b00000000000001100000011111111011;
    assign rom[2821]= 32'b00000000000001100000100111111011;
    assign rom[2822]= 32'b00000000000001100000101111111011;
    assign rom[2823]= 32'b00000000000001100000110111111011;
    assign rom[2824]= 32'b00000000000001100000111111111011;
    assign rom[2825]= 32'b00000000000001100001000111111011;
    assign rom[2826]= 32'b00000000000001100001001111111011;
    assign rom[2827]= 32'b00000000000001100001010111111011;
    assign rom[2828]= 32'b00000000000001100001011111111011;
    assign rom[2829]= 32'b00000000000001100001100111111100;
    assign rom[2830]= 32'b00000000000001100001101111111100;
    assign rom[2831]= 32'b00000000000001100001110111111100;
    assign rom[2832]= 32'b00000000000001100001111111111100;
    assign rom[2833]= 32'b00000000000001100010000111111100;
    assign rom[2834]= 32'b00000000000001100010001111111100;
    assign rom[2835]= 32'b00000000000001100010010111111100;
    assign rom[2836]= 32'b00000000000001100010011111111100;
    assign rom[2837]= 32'b00000000000001100010100111111100;
    assign rom[2838]= 32'b00000000000001100010101111111100;
    assign rom[2839]= 32'b00000000000001100010110111111100;
    assign rom[2840]= 32'b00000000000001100010111111111100;
    assign rom[2841]= 32'b00000000000001100011000111111100;
    assign rom[2842]= 32'b00000000000001100011001111111100;
    assign rom[2843]= 32'b00000000000001100011010111111100;
    assign rom[2844]= 32'b00000000000001100011011111111100;
    assign rom[2845]= 32'b00000000000001100011100111111100;
    assign rom[2846]= 32'b00000000000001100011101111111100;
    assign rom[2847]= 32'b00000000000001100011110111111100;
    assign rom[2848]= 32'b00000000000001100011111111111100;
    assign rom[2849]= 32'b00000000000001100100000111111101;
    assign rom[2850]= 32'b00000000000001100100001111111101;
    assign rom[2851]= 32'b00000000000001100100010111111101;
    assign rom[2852]= 32'b00000000000001100100011111111101;
    assign rom[2853]= 32'b00000000000001100100100111111101;
    assign rom[2854]= 32'b00000000000001100100101111111101;
    assign rom[2855]= 32'b00000000000001100100110111111101;
    assign rom[2856]= 32'b00000000000001100100111111111101;
    assign rom[2857]= 32'b00000000000001100101000111111101;
    assign rom[2858]= 32'b00000000000001100101001111111101;
    assign rom[2859]= 32'b00000000000001100101010111111101;
    assign rom[2860]= 32'b00000000000001100101011111111101;
    assign rom[2861]= 32'b00000000000001100101100111111101;
    assign rom[2862]= 32'b00000000000001100101101111111101;
    assign rom[2863]= 32'b00000000000001100101110111111101;
    assign rom[2864]= 32'b00000000000001100101111111111101;
    assign rom[2865]= 32'b00000000000001100110000111111101;
    assign rom[2866]= 32'b00000000000001100110001111111101;
    assign rom[2867]= 32'b00000000000001100110010111111101;
    assign rom[2868]= 32'b00000000000001100110011111111101;
    assign rom[2869]= 32'b00000000000001100110100111111101;
    assign rom[2870]= 32'b00000000000001100110101111111101;
    assign rom[2871]= 32'b00000000000001100110110111111101;
    assign rom[2872]= 32'b00000000000001100110111111111101;
    assign rom[2873]= 32'b00000000000001100111000111111101;
    assign rom[2874]= 32'b00000000000001100111001111111101;
    assign rom[2875]= 32'b00000000000001100111010111111101;
    assign rom[2876]= 32'b00000000000001100111011111111101;
    assign rom[2877]= 32'b00000000000001100111100111111101;
    assign rom[2878]= 32'b00000000000001100111101111111110;
    assign rom[2879]= 32'b00000000000001100111110111111110;
    assign rom[2880]= 32'b00000000000001100111111111111110;
    assign rom[2881]= 32'b00000000000001101000000111111110;
    assign rom[2882]= 32'b00000000000001101000001111111110;
    assign rom[2883]= 32'b00000000000001101000010111111110;
    assign rom[2884]= 32'b00000000000001101000011111111110;
    assign rom[2885]= 32'b00000000000001101000100111111110;
    assign rom[2886]= 32'b00000000000001101000101111111110;
    assign rom[2887]= 32'b00000000000001101000110111111110;
    assign rom[2888]= 32'b00000000000001101000111111111110;
    assign rom[2889]= 32'b00000000000001101001000111111110;
    assign rom[2890]= 32'b00000000000001101001001111111110;
    assign rom[2891]= 32'b00000000000001101001010111111110;
    assign rom[2892]= 32'b00000000000001101001011111111110;
    assign rom[2893]= 32'b00000000000001101001100111111110;
    assign rom[2894]= 32'b00000000000001101001101111111110;
    assign rom[2895]= 32'b00000000000001101001110111111110;
    assign rom[2896]= 32'b00000000000001101001111111111110;
    assign rom[2897]= 32'b00000000000001101010000111111110;
    assign rom[2898]= 32'b00000000000001101010001111111110;
    assign rom[2899]= 32'b00000000000001101010010111111110;
    assign rom[2900]= 32'b00000000000001101010011111111110;
    assign rom[2901]= 32'b00000000000001101010100111111110;
    assign rom[2902]= 32'b00000000000001101010101111111110;
    assign rom[2903]= 32'b00000000000001101010110111111110;
    assign rom[2904]= 32'b00000000000001101010111111111110;
    assign rom[2905]= 32'b00000000000001101011000111111110;
    assign rom[2906]= 32'b00000000000001101011001111111110;
    assign rom[2907]= 32'b00000000000001101011010111111110;
    assign rom[2908]= 32'b00000000000001101011011111111110;
    assign rom[2909]= 32'b00000000000001101011100111111110;
    assign rom[2910]= 32'b00000000000001101011101111111110;
    assign rom[2911]= 32'b00000000000001101011110111111110;
    assign rom[2912]= 32'b00000000000001101011111111111110;
    assign rom[2913]= 32'b00000000000001101100000111111110;
    assign rom[2914]= 32'b00000000000001101100001111111110;
    assign rom[2915]= 32'b00000000000001101100010111111110;
    assign rom[2916]= 32'b00000000000001101100011111111110;
    assign rom[2917]= 32'b00000000000001101100100111111110;
    assign rom[2918]= 32'b00000000000001101100101111111110;
    assign rom[2919]= 32'b00000000000001101100110111111110;
    assign rom[2920]= 32'b00000000000001101100111111111110;
    assign rom[2921]= 32'b00000000000001101101000111111110;
    assign rom[2922]= 32'b00000000000001101101001111111110;
    assign rom[2923]= 32'b00000000000001101101010111111110;
    assign rom[2924]= 32'b00000000000001101101011111111110;
    assign rom[2925]= 32'b00000000000001101101100111111110;
    assign rom[2926]= 32'b00000000000001101101101111111111;
    assign rom[2927]= 32'b00000000000001101101110111111111;
    assign rom[2928]= 32'b00000000000001101101111111111111;
    assign rom[2929]= 32'b00000000000001101110000111111111;
    assign rom[2930]= 32'b00000000000001101110001111111111;
    assign rom[2931]= 32'b00000000000001101110010111111111;
    assign rom[2932]= 32'b00000000000001101110011111111111;
    assign rom[2933]= 32'b00000000000001101110100111111111;
    assign rom[2934]= 32'b00000000000001101110101111111111;
    assign rom[2935]= 32'b00000000000001101110110111111111;
    assign rom[2936]= 32'b00000000000001101110111111111111;
    assign rom[2937]= 32'b00000000000001101111000111111111;
    assign rom[2938]= 32'b00000000000001101111001111111111;
    assign rom[2939]= 32'b00000000000001101111010111111111;
    assign rom[2940]= 32'b00000000000001101111011111111111;
    assign rom[2941]= 32'b00000000000001101111100111111111;
    assign rom[2942]= 32'b00000000000001101111101111111111;
    assign rom[2943]= 32'b00000000000001101111110111111111;
    assign rom[2944]= 32'b00000000000001101111111111111111;
    assign rom[2945]= 32'b00000000000001110000000111111111;
    assign rom[2946]= 32'b00000000000001110000001111111111;
    assign rom[2947]= 32'b00000000000001110000010111111111;
    assign rom[2948]= 32'b00000000000001110000011111111111;
    assign rom[2949]= 32'b00000000000001110000100111111111;
    assign rom[2950]= 32'b00000000000001110000101111111111;
    assign rom[2951]= 32'b00000000000001110000110111111111;
    assign rom[2952]= 32'b00000000000001110000111111111111;
    assign rom[2953]= 32'b00000000000001110001000111111111;
    assign rom[2954]= 32'b00000000000001110001001111111111;
    assign rom[2955]= 32'b00000000000001110001010111111111;
    assign rom[2956]= 32'b00000000000001110001011111111111;
    assign rom[2957]= 32'b00000000000001110001100111111111;
    assign rom[2958]= 32'b00000000000001110001101111111111;
    assign rom[2959]= 32'b00000000000001110001110111111111;
    assign rom[2960]= 32'b00000000000001110001111111111111;
    assign rom[2961]= 32'b00000000000001110010000111111111;
    assign rom[2962]= 32'b00000000000001110010001111111111;
    assign rom[2963]= 32'b00000000000001110010010111111111;
    assign rom[2964]= 32'b00000000000001110010011111111111;
    assign rom[2965]= 32'b00000000000001110010100111111111;
    assign rom[2966]= 32'b00000000000001110010101111111111;
    assign rom[2967]= 32'b00000000000001110010110111111111;
    assign rom[2968]= 32'b00000000000001110010111111111111;
    assign rom[2969]= 32'b00000000000001110011000111111111;
    assign rom[2970]= 32'b00000000000001110011001111111111;
    assign rom[2971]= 32'b00000000000001110011010111111111;
    assign rom[2972]= 32'b00000000000001110011011111111111;
    assign rom[2973]= 32'b00000000000001110011100111111111;
    assign rom[2974]= 32'b00000000000001110011101111111111;
    assign rom[2975]= 32'b00000000000001110011110111111111;
    assign rom[2976]= 32'b00000000000001110011111111111111;
    assign rom[2977]= 32'b00000000000001110100000111111111;
    assign rom[2978]= 32'b00000000000001110100001111111111;
    assign rom[2979]= 32'b00000000000001110100010111111111;
    assign rom[2980]= 32'b00000000000001110100011111111111;
    assign rom[2981]= 32'b00000000000001110100100111111111;
    assign rom[2982]= 32'b00000000000001110100101111111111;
    assign rom[2983]= 32'b00000000000001110100110111111111;
    assign rom[2984]= 32'b00000000000001110100111111111111;
    assign rom[2985]= 32'b00000000000001110101000111111111;
    assign rom[2986]= 32'b00000000000001110101001111111111;
    assign rom[2987]= 32'b00000000000001110101010111111111;
    assign rom[2988]= 32'b00000000000001110101011111111111;
    assign rom[2989]= 32'b00000000000001110101100111111111;
    assign rom[2990]= 32'b00000000000001110101101111111111;
    assign rom[2991]= 32'b00000000000001110101110111111111;
    assign rom[2992]= 32'b00000000000001110101111111111111;
    assign rom[2993]= 32'b00000000000001110110000111111111;
    assign rom[2994]= 32'b00000000000001110110001111111111;
    assign rom[2995]= 32'b00000000000001110110010111111111;
    assign rom[2996]= 32'b00000000000001110110011111111111;
    assign rom[2997]= 32'b00000000000001110110100111111111;
    assign rom[2998]= 32'b00000000000001110110101111111111;
    assign rom[2999]= 32'b00000000000001110110110111111111;
    assign rom[3000]= 32'b00000000000001110110111111111111;
    assign rom[3001]= 32'b00000000000001110111000111111111;
    assign rom[3002]= 32'b00000000000001110111001111111111;
    assign rom[3003]= 32'b00000000000001110111010111111111;
    assign rom[3004]= 32'b00000000000001110111011111111111;
    assign rom[3005]= 32'b00000000000001110111100111111111;
    assign rom[3006]= 32'b00000000000001110111101111111111;
    assign rom[3007]= 32'b00000000000001110111110111111111;
    assign rom[3008]= 32'b00000000000001110111111111111111;
    assign rom[3009]= 32'b00000000000001111000000111111111;
    assign rom[3010]= 32'b00000000000001111000001111111111;
    assign rom[3011]= 32'b00000000000001111000010111111111;
    assign rom[3012]= 32'b00000000000001111000011111111111;
    assign rom[3013]= 32'b00000000000001111000100111111111;
    assign rom[3014]= 32'b00000000000001111000101111111111;
    assign rom[3015]= 32'b00000000000001111000110111111111;
    assign rom[3016]= 32'b00000000000001111000111111111111;
    assign rom[3017]= 32'b00000000000001111001000111111111;
    assign rom[3018]= 32'b00000000000001111001001111111111;
    assign rom[3019]= 32'b00000000000001111001010111111111;
    assign rom[3020]= 32'b00000000000001111001011111111111;
    assign rom[3021]= 32'b00000000000001111001100111111111;
    assign rom[3022]= 32'b00000000000001111001101111111111;
    assign rom[3023]= 32'b00000000000001111001110111111111;
    assign rom[3024]= 32'b00000000000001111001111111111111;
    assign rom[3025]= 32'b00000000000001111010000111111111;
    assign rom[3026]= 32'b00000000000001111010001111111111;
    assign rom[3027]= 32'b00000000000001111010010111111111;
    assign rom[3028]= 32'b00000000000001111010011111111111;
    assign rom[3029]= 32'b00000000000001111010100111111111;
    assign rom[3030]= 32'b00000000000001111010101111111111;
    assign rom[3031]= 32'b00000000000001111010110111111111;
    assign rom[3032]= 32'b00000000000001111010111111111111;
    assign rom[3033]= 32'b00000000000001111011000111111111;
    assign rom[3034]= 32'b00000000000001111011001111111111;
    assign rom[3035]= 32'b00000000000001111011010111111111;
    assign rom[3036]= 32'b00000000000001111011011111111111;
    assign rom[3037]= 32'b00000000000001111011100111111111;
    assign rom[3038]= 32'b00000000000001111011101111111111;
    assign rom[3039]= 32'b00000000000001111011110111111111;
    assign rom[3040]= 32'b00000000000001111011111111111111;
    assign rom[3041]= 32'b00000000000001111100000111111111;
    assign rom[3042]= 32'b00000000000001111100001111111111;
    assign rom[3043]= 32'b00000000000001111100010111111111;
    assign rom[3044]= 32'b00000000000001111100011111111111;
    assign rom[3045]= 32'b00000000000001111100100111111111;
    assign rom[3046]= 32'b00000000000001111100101111111111;
    assign rom[3047]= 32'b00000000000001111100110111111111;
    assign rom[3048]= 32'b00000000000001111100111111111111;
    assign rom[3049]= 32'b00000000000001111101000111111111;
    assign rom[3050]= 32'b00000000000001111101001111111111;
    assign rom[3051]= 32'b00000000000001111101010111111111;
    assign rom[3052]= 32'b00000000000001111101011111111111;
    assign rom[3053]= 32'b00000000000001111101100111111111;
    assign rom[3054]= 32'b00000000000001111101101111111111;
    assign rom[3055]= 32'b00000000000001111101110111111111;
    assign rom[3056]= 32'b00000000000001111101111111111111;
    assign rom[3057]= 32'b00000000000001111110000111111111;
    assign rom[3058]= 32'b00000000000001111110001111111111;
    assign rom[3059]= 32'b00000000000001111110010111111111;
    assign rom[3060]= 32'b00000000000001111110011111111111;
    assign rom[3061]= 32'b00000000000001111110100111111111;
    assign rom[3062]= 32'b00000000000001111110101111111111;
    assign rom[3063]= 32'b00000000000001111110110111111111;
    assign rom[3064]= 32'b00000000000001111110111111111111;
    assign rom[3065]= 32'b00000000000001111111000111111111;
    assign rom[3066]= 32'b00000000000001111111001111111111;
    assign rom[3067]= 32'b00000000000001111111010111111111;
    assign rom[3068]= 32'b00000000000001111111011111111111;
    assign rom[3069]= 32'b00000000000001111111100111111111;
    assign rom[3070]= 32'b00000000000001111111101111111111;
    assign rom[3071]= 32'b00000000000001111111110111111111;
    assign rom[3072]= 32'b00000000000001111111111111111111;
    assign rom[3073]= 32'b00000000000010000000000111111111;
    assign rom[3074]= 32'b00000000000010000000001111111111;
    assign rom[3075]= 32'b00000000000010000000010111111111;
    assign rom[3076]= 32'b00000000000010000000011111111111;
    assign rom[3077]= 32'b00000000000010000000100111111111;
    assign rom[3078]= 32'b00000000000010000000101111111111;
    assign rom[3079]= 32'b00000000000010000000110111111111;
    assign rom[3080]= 32'b00000000000010000000111111111111;
    assign rom[3081]= 32'b00000000000010000001000111111111;
    assign rom[3082]= 32'b00000000000010000001001111111111;
    assign rom[3083]= 32'b00000000000010000001010111111111;
    assign rom[3084]= 32'b00000000000010000001011111111111;
    assign rom[3085]= 32'b00000000000010000001100111111111;
    assign rom[3086]= 32'b00000000000010000001101111111111;
    assign rom[3087]= 32'b00000000000010000001110111111111;
    assign rom[3088]= 32'b00000000000010000001111111111111;
    assign rom[3089]= 32'b00000000000010000010000111111111;
    assign rom[3090]= 32'b00000000000010000010001111111111;
    assign rom[3091]= 32'b00000000000010000010010111111111;
    assign rom[3092]= 32'b00000000000010000010011111111111;
    assign rom[3093]= 32'b00000000000010000010100111111111;
    assign rom[3094]= 32'b00000000000010000010101111111111;
    assign rom[3095]= 32'b00000000000010000010110111111111;
    assign rom[3096]= 32'b00000000000010000010111111111111;
    assign rom[3097]= 32'b00000000000010000011000111111111;
    assign rom[3098]= 32'b00000000000010000011001111111111;
    assign rom[3099]= 32'b00000000000010000011010111111111;
    assign rom[3100]= 32'b00000000000010000011011111111111;
    assign rom[3101]= 32'b00000000000010000011100111111111;
    assign rom[3102]= 32'b00000000000010000011101111111111;
    assign rom[3103]= 32'b00000000000010000011110111111111;
    assign rom[3104]= 32'b00000000000010000011111111111111;
    assign rom[3105]= 32'b00000000000010000100000111111111;
    assign rom[3106]= 32'b00000000000010000100001111111111;
    assign rom[3107]= 32'b00000000000010000100010111111111;
    assign rom[3108]= 32'b00000000000010000100011111111111;
    assign rom[3109]= 32'b00000000000010000100100111111111;
    assign rom[3110]= 32'b00000000000010000100101111111111;
    assign rom[3111]= 32'b00000000000010000100110111111111;
    assign rom[3112]= 32'b00000000000010000100111111111111;
    assign rom[3113]= 32'b00000000000010000101000111111111;
    assign rom[3114]= 32'b00000000000010000101001111111111;
    assign rom[3115]= 32'b00000000000010000101010111111111;
    assign rom[3116]= 32'b00000000000010000101011111111111;
    assign rom[3117]= 32'b00000000000010000101100111111111;
    assign rom[3118]= 32'b00000000000010000101101111111111;
    assign rom[3119]= 32'b00000000000010000101110111111111;
    assign rom[3120]= 32'b00000000000010000101111111111111;
    assign rom[3121]= 32'b00000000000010000110000111111111;
    assign rom[3122]= 32'b00000000000010000110001111111111;
    assign rom[3123]= 32'b00000000000010000110010111111111;
    assign rom[3124]= 32'b00000000000010000110011111111111;
    assign rom[3125]= 32'b00000000000010000110100111111111;
    assign rom[3126]= 32'b00000000000010000110101111111111;
    assign rom[3127]= 32'b00000000000010000110110111111111;
    assign rom[3128]= 32'b00000000000010000110111111111111;
    assign rom[3129]= 32'b00000000000010000111000111111111;
    assign rom[3130]= 32'b00000000000010000111001111111111;
    assign rom[3131]= 32'b00000000000010000111010111111111;
    assign rom[3132]= 32'b00000000000010000111011111111111;
    assign rom[3133]= 32'b00000000000010000111100111111111;
    assign rom[3134]= 32'b00000000000010000111101111111111;
    assign rom[3135]= 32'b00000000000010000111110111111111;
    assign rom[3136]= 32'b00000000000010000111111111111111;
    assign rom[3137]= 32'b00000000000010001000000111111111;
    assign rom[3138]= 32'b00000000000010001000001111111111;
    assign rom[3139]= 32'b00000000000010001000010111111111;
    assign rom[3140]= 32'b00000000000010001000011111111111;
    assign rom[3141]= 32'b00000000000010001000100111111111;
    assign rom[3142]= 32'b00000000000010001000101111111111;
    assign rom[3143]= 32'b00000000000010001000110111111111;
    assign rom[3144]= 32'b00000000000010001000111111111111;
    assign rom[3145]= 32'b00000000000010001001000111111111;
    assign rom[3146]= 32'b00000000000010001001001111111111;
    assign rom[3147]= 32'b00000000000010001001010111111111;
    assign rom[3148]= 32'b00000000000010001001011111111111;
    assign rom[3149]= 32'b00000000000010001001100111111111;
    assign rom[3150]= 32'b00000000000010001001101111111111;
    assign rom[3151]= 32'b00000000000010001001110111111111;
    assign rom[3152]= 32'b00000000000010001001111111111111;
    assign rom[3153]= 32'b00000000000010001010000111111111;
    assign rom[3154]= 32'b00000000000010001010001111111111;
    assign rom[3155]= 32'b00000000000010001010010111111111;
    assign rom[3156]= 32'b00000000000010001010011111111111;
    assign rom[3157]= 32'b00000000000010001010100111111111;
    assign rom[3158]= 32'b00000000000010001010101111111111;
    assign rom[3159]= 32'b00000000000010001010110111111111;
    assign rom[3160]= 32'b00000000000010001010111111111111;
    assign rom[3161]= 32'b00000000000010001011000111111111;
    assign rom[3162]= 32'b00000000000010001011001111111111;
    assign rom[3163]= 32'b00000000000010001011010111111111;
    assign rom[3164]= 32'b00000000000010001011011111111111;
    assign rom[3165]= 32'b00000000000010001011100111111111;
    assign rom[3166]= 32'b00000000000010001011101111111111;
    assign rom[3167]= 32'b00000000000010001011110111111111;
    assign rom[3168]= 32'b00000000000010001011111111111111;
    assign rom[3169]= 32'b00000000000010001100000111111111;
    assign rom[3170]= 32'b00000000000010001100001111111111;
    assign rom[3171]= 32'b00000000000010001100010111111111;
    assign rom[3172]= 32'b00000000000010001100011111111111;
    assign rom[3173]= 32'b00000000000010001100100111111111;
    assign rom[3174]= 32'b00000000000010001100101111111111;
    assign rom[3175]= 32'b00000000000010001100110111111111;
    assign rom[3176]= 32'b00000000000010001100111111111111;
    assign rom[3177]= 32'b00000000000010001101000111111111;
    assign rom[3178]= 32'b00000000000010001101001111111111;
    assign rom[3179]= 32'b00000000000010001101010111111111;
    assign rom[3180]= 32'b00000000000010001101011111111111;
    assign rom[3181]= 32'b00000000000010001101100111111111;
    assign rom[3182]= 32'b00000000000010001101101111111111;
    assign rom[3183]= 32'b00000000000010001101110111111111;
    assign rom[3184]= 32'b00000000000010001101111111111111;
    assign rom[3185]= 32'b00000000000010001110000111111111;
    assign rom[3186]= 32'b00000000000010001110001111111111;
    assign rom[3187]= 32'b00000000000010001110010111111111;
    assign rom[3188]= 32'b00000000000010001110011111111111;
    assign rom[3189]= 32'b00000000000010001110100111111111;
    assign rom[3190]= 32'b00000000000010001110101111111111;
    assign rom[3191]= 32'b00000000000010001110110111111111;
    assign rom[3192]= 32'b00000000000010001110111111111111;
    assign rom[3193]= 32'b00000000000010001111000111111111;
    assign rom[3194]= 32'b00000000000010001111001111111111;
    assign rom[3195]= 32'b00000000000010001111010111111111;
    assign rom[3196]= 32'b00000000000010001111011111111111;
    assign rom[3197]= 32'b00000000000010001111100111111111;
    assign rom[3198]= 32'b00000000000010001111101111111111;
    assign rom[3199]= 32'b00000000000010001111110111111111;
    assign rom[3200]= 32'b00000000000010001111111111111111;
    assign rom[3201]= 32'b00000000000010010000000111111111;
    assign rom[3202]= 32'b00000000000010010000001111111111;
    assign rom[3203]= 32'b00000000000010010000010111111111;
    assign rom[3204]= 32'b00000000000010010000011111111111;
    assign rom[3205]= 32'b00000000000010010000100111111111;
    assign rom[3206]= 32'b00000000000010010000101111111111;
    assign rom[3207]= 32'b00000000000010010000110111111111;
    assign rom[3208]= 32'b00000000000010010000111111111111;
    assign rom[3209]= 32'b00000000000010010001000111111111;
    assign rom[3210]= 32'b00000000000010010001001111111111;
    assign rom[3211]= 32'b00000000000010010001010111111111;
    assign rom[3212]= 32'b00000000000010010001011111111111;
    assign rom[3213]= 32'b00000000000010010001100111111111;
    assign rom[3214]= 32'b00000000000010010001101111111111;
    assign rom[3215]= 32'b00000000000010010001110111111111;
    assign rom[3216]= 32'b00000000000010010001111111111111;
    assign rom[3217]= 32'b00000000000010010010000111111111;
    assign rom[3218]= 32'b00000000000010010010001111111111;
    assign rom[3219]= 32'b00000000000010010010010111111111;
    assign rom[3220]= 32'b00000000000010010010011111111111;
    assign rom[3221]= 32'b00000000000010010010100111111111;
    assign rom[3222]= 32'b00000000000010010010101111111111;
    assign rom[3223]= 32'b00000000000010010010110111111111;
    assign rom[3224]= 32'b00000000000010010010111111111111;
    assign rom[3225]= 32'b00000000000010010011000111111111;
    assign rom[3226]= 32'b00000000000010010011001111111111;
    assign rom[3227]= 32'b00000000000010010011010111111111;
    assign rom[3228]= 32'b00000000000010010011011111111111;
    assign rom[3229]= 32'b00000000000010010011100111111111;
    assign rom[3230]= 32'b00000000000010010011101111111111;
    assign rom[3231]= 32'b00000000000010010011110111111111;
    assign rom[3232]= 32'b00000000000010010011111111111111;
    assign rom[3233]= 32'b00000000000010010100000111111111;
    assign rom[3234]= 32'b00000000000010010100001111111111;
    assign rom[3235]= 32'b00000000000010010100010111111111;
    assign rom[3236]= 32'b00000000000010010100011111111111;
    assign rom[3237]= 32'b00000000000010010100100111111111;
    assign rom[3238]= 32'b00000000000010010100101111111111;
    assign rom[3239]= 32'b00000000000010010100110111111111;
    assign rom[3240]= 32'b00000000000010010100111111111111;
    assign rom[3241]= 32'b00000000000010010101000111111111;
    assign rom[3242]= 32'b00000000000010010101001111111111;
    assign rom[3243]= 32'b00000000000010010101010111111111;
    assign rom[3244]= 32'b00000000000010010101011111111111;
    assign rom[3245]= 32'b00000000000010010101100111111111;
    assign rom[3246]= 32'b00000000000010010101101111111111;
    assign rom[3247]= 32'b00000000000010010101110111111111;
    assign rom[3248]= 32'b00000000000010010101111111111111;
    assign rom[3249]= 32'b00000000000010010110000111111111;
    assign rom[3250]= 32'b00000000000010010110001111111111;
    assign rom[3251]= 32'b00000000000010010110010111111111;
    assign rom[3252]= 32'b00000000000010010110011111111111;
    assign rom[3253]= 32'b00000000000010010110100111111111;
    assign rom[3254]= 32'b00000000000010010110101111111111;
    assign rom[3255]= 32'b00000000000010010110110111111111;
    assign rom[3256]= 32'b00000000000010010110111111111111;
    assign rom[3257]= 32'b00000000000010010111000111111111;
    assign rom[3258]= 32'b00000000000010010111001111111111;
    assign rom[3259]= 32'b00000000000010010111010111111111;
    assign rom[3260]= 32'b00000000000010010111011111111111;
    assign rom[3261]= 32'b00000000000010010111100111111111;
    assign rom[3262]= 32'b00000000000010010111101111111111;
    assign rom[3263]= 32'b00000000000010010111110111111111;
    assign rom[3264]= 32'b00000000000010010111111111111111;
    assign rom[3265]= 32'b00000000000010011000000111111111;
    assign rom[3266]= 32'b00000000000010011000001111111111;
    assign rom[3267]= 32'b00000000000010011000010111111111;
    assign rom[3268]= 32'b00000000000010011000011111111111;
    assign rom[3269]= 32'b00000000000010011000100111111111;
    assign rom[3270]= 32'b00000000000010011000101111111111;
    assign rom[3271]= 32'b00000000000010011000110111111111;
    assign rom[3272]= 32'b00000000000010011000111111111111;
    assign rom[3273]= 32'b00000000000010011001000111111111;
    assign rom[3274]= 32'b00000000000010011001001111111111;
    assign rom[3275]= 32'b00000000000010011001010111111111;
    assign rom[3276]= 32'b00000000000010011001011111111111;
    assign rom[3277]= 32'b00000000000010011001100111111111;
    assign rom[3278]= 32'b00000000000010011001101111111111;
    assign rom[3279]= 32'b00000000000010011001110111111111;
    assign rom[3280]= 32'b00000000000010011001111111111111;
    assign rom[3281]= 32'b00000000000010011010000111111111;
    assign rom[3282]= 32'b00000000000010011010001111111111;
    assign rom[3283]= 32'b00000000000010011010010111111111;
    assign rom[3284]= 32'b00000000000010011010011111111111;
    assign rom[3285]= 32'b00000000000010011010100111111111;
    assign rom[3286]= 32'b00000000000010011010101111111111;
    assign rom[3287]= 32'b00000000000010011010110111111111;
    assign rom[3288]= 32'b00000000000010011010111111111111;
    assign rom[3289]= 32'b00000000000010011011000111111111;
    assign rom[3290]= 32'b00000000000010011011001111111111;
    assign rom[3291]= 32'b00000000000010011011010111111111;
    assign rom[3292]= 32'b00000000000010011011011111111111;
    assign rom[3293]= 32'b00000000000010011011100111111111;
    assign rom[3294]= 32'b00000000000010011011101111111111;
    assign rom[3295]= 32'b00000000000010011011110111111111;
    assign rom[3296]= 32'b00000000000010011011111111111111;
    assign rom[3297]= 32'b00000000000010011100000111111111;
    assign rom[3298]= 32'b00000000000010011100001111111111;
    assign rom[3299]= 32'b00000000000010011100010111111111;
    assign rom[3300]= 32'b00000000000010011100011111111111;
    assign rom[3301]= 32'b00000000000010011100100111111111;
    assign rom[3302]= 32'b00000000000010011100101111111111;
    assign rom[3303]= 32'b00000000000010011100110111111111;
    assign rom[3304]= 32'b00000000000010011100111111111111;
    assign rom[3305]= 32'b00000000000010011101000111111111;
    assign rom[3306]= 32'b00000000000010011101001111111111;
    assign rom[3307]= 32'b00000000000010011101010111111111;
    assign rom[3308]= 32'b00000000000010011101011111111111;
    assign rom[3309]= 32'b00000000000010011101100111111111;
    assign rom[3310]= 32'b00000000000010011101101111111111;
    assign rom[3311]= 32'b00000000000010011101110111111111;
    assign rom[3312]= 32'b00000000000010011101111111111111;
    assign rom[3313]= 32'b00000000000010011110000111111111;
    assign rom[3314]= 32'b00000000000010011110001111111111;
    assign rom[3315]= 32'b00000000000010011110010111111111;
    assign rom[3316]= 32'b00000000000010011110011111111111;
    assign rom[3317]= 32'b00000000000010011110100111111111;
    assign rom[3318]= 32'b00000000000010011110101111111111;
    assign rom[3319]= 32'b00000000000010011110110111111111;
    assign rom[3320]= 32'b00000000000010011110111111111111;
    assign rom[3321]= 32'b00000000000010011111000111111111;
    assign rom[3322]= 32'b00000000000010011111001111111111;
    assign rom[3323]= 32'b00000000000010011111010111111111;
    assign rom[3324]= 32'b00000000000010011111011111111111;
    assign rom[3325]= 32'b00000000000010011111100111111111;
    assign rom[3326]= 32'b00000000000010011111101111111111;
    assign rom[3327]= 32'b00000000000010011111110111111111;
    assign rom[3328]= 32'b00000000000010011111111111111111;
    assign rom[3329]= 32'b00000000000010100000000111111111;
    assign rom[3330]= 32'b00000000000010100000001111111111;
    assign rom[3331]= 32'b00000000000010100000010111111111;
    assign rom[3332]= 32'b00000000000010100000011111111111;
    assign rom[3333]= 32'b00000000000010100000100111111111;
    assign rom[3334]= 32'b00000000000010100000101111111111;
    assign rom[3335]= 32'b00000000000010100000110111111111;
    assign rom[3336]= 32'b00000000000010100000111111111111;
    assign rom[3337]= 32'b00000000000010100001000111111111;
    assign rom[3338]= 32'b00000000000010100001001111111111;
    assign rom[3339]= 32'b00000000000010100001010111111111;
    assign rom[3340]= 32'b00000000000010100001011111111111;
    assign rom[3341]= 32'b00000000000010100001100111111111;
    assign rom[3342]= 32'b00000000000010100001101111111111;
    assign rom[3343]= 32'b00000000000010100001110111111111;
    assign rom[3344]= 32'b00000000000010100001111111111111;
    assign rom[3345]= 32'b00000000000010100010000111111111;
    assign rom[3346]= 32'b00000000000010100010001111111111;
    assign rom[3347]= 32'b00000000000010100010010111111111;
    assign rom[3348]= 32'b00000000000010100010011111111111;
    assign rom[3349]= 32'b00000000000010100010100111111111;
    assign rom[3350]= 32'b00000000000010100010101111111111;
    assign rom[3351]= 32'b00000000000010100010110111111111;
    assign rom[3352]= 32'b00000000000010100010111111111111;
    assign rom[3353]= 32'b00000000000010100011000111111111;
    assign rom[3354]= 32'b00000000000010100011001111111111;
    assign rom[3355]= 32'b00000000000010100011010111111111;
    assign rom[3356]= 32'b00000000000010100011011111111111;
    assign rom[3357]= 32'b00000000000010100011100111111111;
    assign rom[3358]= 32'b00000000000010100011101111111111;
    assign rom[3359]= 32'b00000000000010100011110111111111;
    assign rom[3360]= 32'b00000000000010100011111111111111;
    assign rom[3361]= 32'b00000000000010100100000111111111;
    assign rom[3362]= 32'b00000000000010100100001111111111;
    assign rom[3363]= 32'b00000000000010100100010111111111;
    assign rom[3364]= 32'b00000000000010100100011111111111;
    assign rom[3365]= 32'b00000000000010100100100111111111;
    assign rom[3366]= 32'b00000000000010100100101111111111;
    assign rom[3367]= 32'b00000000000010100100110111111111;
    assign rom[3368]= 32'b00000000000010100100111111111111;
    assign rom[3369]= 32'b00000000000010100101000111111111;
    assign rom[3370]= 32'b00000000000010100101001111111111;
    assign rom[3371]= 32'b00000000000010100101010111111111;
    assign rom[3372]= 32'b00000000000010100101011111111111;
    assign rom[3373]= 32'b00000000000010100101100111111111;
    assign rom[3374]= 32'b00000000000010100101101111111111;
    assign rom[3375]= 32'b00000000000010100101110111111111;
    assign rom[3376]= 32'b00000000000010100101111111111111;
    assign rom[3377]= 32'b00000000000010100110000111111111;
    assign rom[3378]= 32'b00000000000010100110001111111111;
    assign rom[3379]= 32'b00000000000010100110010111111111;
    assign rom[3380]= 32'b00000000000010100110011111111111;
    assign rom[3381]= 32'b00000000000010100110100111111111;
    assign rom[3382]= 32'b00000000000010100110101111111111;
    assign rom[3383]= 32'b00000000000010100110110111111111;
    assign rom[3384]= 32'b00000000000010100110111111111111;
    assign rom[3385]= 32'b00000000000010100111000111111111;
    assign rom[3386]= 32'b00000000000010100111001111111111;
    assign rom[3387]= 32'b00000000000010100111010111111111;
    assign rom[3388]= 32'b00000000000010100111011111111111;
    assign rom[3389]= 32'b00000000000010100111100111111111;
    assign rom[3390]= 32'b00000000000010100111101111111111;
    assign rom[3391]= 32'b00000000000010100111110111111111;
    assign rom[3392]= 32'b00000000000010100111111111111111;
    assign rom[3393]= 32'b00000000000010101000000111111111;
    assign rom[3394]= 32'b00000000000010101000001111111111;
    assign rom[3395]= 32'b00000000000010101000010111111111;
    assign rom[3396]= 32'b00000000000010101000011111111111;
    assign rom[3397]= 32'b00000000000010101000100111111111;
    assign rom[3398]= 32'b00000000000010101000101111111111;
    assign rom[3399]= 32'b00000000000010101000110111111111;
    assign rom[3400]= 32'b00000000000010101000111111111111;
    assign rom[3401]= 32'b00000000000010101001000111111111;
    assign rom[3402]= 32'b00000000000010101001001111111111;
    assign rom[3403]= 32'b00000000000010101001010111111111;
    assign rom[3404]= 32'b00000000000010101001011111111111;
    assign rom[3405]= 32'b00000000000010101001100111111111;
    assign rom[3406]= 32'b00000000000010101001101111111111;
    assign rom[3407]= 32'b00000000000010101001110111111111;
    assign rom[3408]= 32'b00000000000010101001111111111111;
    assign rom[3409]= 32'b00000000000010101010000111111111;
    assign rom[3410]= 32'b00000000000010101010001111111111;
    assign rom[3411]= 32'b00000000000010101010010111111111;
    assign rom[3412]= 32'b00000000000010101010011111111111;
    assign rom[3413]= 32'b00000000000010101010100111111111;
    assign rom[3414]= 32'b00000000000010101010101111111111;
    assign rom[3415]= 32'b00000000000010101010110111111111;
    assign rom[3416]= 32'b00000000000010101010111111111111;
    assign rom[3417]= 32'b00000000000010101011000111111111;
    assign rom[3418]= 32'b00000000000010101011001111111111;
    assign rom[3419]= 32'b00000000000010101011010111111111;
    assign rom[3420]= 32'b00000000000010101011011111111111;
    assign rom[3421]= 32'b00000000000010101011100111111111;
    assign rom[3422]= 32'b00000000000010101011101111111111;
    assign rom[3423]= 32'b00000000000010101011110111111111;
    assign rom[3424]= 32'b00000000000010101011111111111111;
    assign rom[3425]= 32'b00000000000010101100000111111111;
    assign rom[3426]= 32'b00000000000010101100001111111111;
    assign rom[3427]= 32'b00000000000010101100010111111111;
    assign rom[3428]= 32'b00000000000010101100011111111111;
    assign rom[3429]= 32'b00000000000010101100100111111111;
    assign rom[3430]= 32'b00000000000010101100101111111111;
    assign rom[3431]= 32'b00000000000010101100110111111111;
    assign rom[3432]= 32'b00000000000010101100111111111111;
    assign rom[3433]= 32'b00000000000010101101000111111111;
    assign rom[3434]= 32'b00000000000010101101001111111111;
    assign rom[3435]= 32'b00000000000010101101010111111111;
    assign rom[3436]= 32'b00000000000010101101011111111111;
    assign rom[3437]= 32'b00000000000010101101100111111111;
    assign rom[3438]= 32'b00000000000010101101101111111111;
    assign rom[3439]= 32'b00000000000010101101110111111111;
    assign rom[3440]= 32'b00000000000010101101111111111111;
    assign rom[3441]= 32'b00000000000010101110000111111111;
    assign rom[3442]= 32'b00000000000010101110001111111111;
    assign rom[3443]= 32'b00000000000010101110010111111111;
    assign rom[3444]= 32'b00000000000010101110011111111111;
    assign rom[3445]= 32'b00000000000010101110100111111111;
    assign rom[3446]= 32'b00000000000010101110101111111111;
    assign rom[3447]= 32'b00000000000010101110110111111111;
    assign rom[3448]= 32'b00000000000010101110111111111111;
    assign rom[3449]= 32'b00000000000010101111000111111111;
    assign rom[3450]= 32'b00000000000010101111001111111111;
    assign rom[3451]= 32'b00000000000010101111010111111111;
    assign rom[3452]= 32'b00000000000010101111011111111111;
    assign rom[3453]= 32'b00000000000010101111100111111111;
    assign rom[3454]= 32'b00000000000010101111101111111111;
    assign rom[3455]= 32'b00000000000010101111110111111111;
    assign rom[3456]= 32'b00000000000010101111111111111111;
    assign rom[3457]= 32'b00000000000010110000000111111111;
    assign rom[3458]= 32'b00000000000010110000001111111111;
    assign rom[3459]= 32'b00000000000010110000010111111111;
    assign rom[3460]= 32'b00000000000010110000011111111111;
    assign rom[3461]= 32'b00000000000010110000100111111111;
    assign rom[3462]= 32'b00000000000010110000101111111111;
    assign rom[3463]= 32'b00000000000010110000110111111111;
    assign rom[3464]= 32'b00000000000010110000111111111111;
    assign rom[3465]= 32'b00000000000010110001000111111111;
    assign rom[3466]= 32'b00000000000010110001001111111111;
    assign rom[3467]= 32'b00000000000010110001010111111111;
    assign rom[3468]= 32'b00000000000010110001011111111111;
    assign rom[3469]= 32'b00000000000010110001100111111111;
    assign rom[3470]= 32'b00000000000010110001101111111111;
    assign rom[3471]= 32'b00000000000010110001110111111111;
    assign rom[3472]= 32'b00000000000010110001111111111111;
    assign rom[3473]= 32'b00000000000010110010000111111111;
    assign rom[3474]= 32'b00000000000010110010001111111111;
    assign rom[3475]= 32'b00000000000010110010010111111111;
    assign rom[3476]= 32'b00000000000010110010011111111111;
    assign rom[3477]= 32'b00000000000010110010100111111111;
    assign rom[3478]= 32'b00000000000010110010101111111111;
    assign rom[3479]= 32'b00000000000010110010110111111111;
    assign rom[3480]= 32'b00000000000010110010111111111111;
    assign rom[3481]= 32'b00000000000010110011000111111111;
    assign rom[3482]= 32'b00000000000010110011001111111111;
    assign rom[3483]= 32'b00000000000010110011010111111111;
    assign rom[3484]= 32'b00000000000010110011011111111111;
    assign rom[3485]= 32'b00000000000010110011100111111111;
    assign rom[3486]= 32'b00000000000010110011101111111111;
    assign rom[3487]= 32'b00000000000010110011110111111111;
    assign rom[3488]= 32'b00000000000010110011111111111111;
    assign rom[3489]= 32'b00000000000010110100000111111111;
    assign rom[3490]= 32'b00000000000010110100001111111111;
    assign rom[3491]= 32'b00000000000010110100010111111111;
    assign rom[3492]= 32'b00000000000010110100011111111111;
    assign rom[3493]= 32'b00000000000010110100100111111111;
    assign rom[3494]= 32'b00000000000010110100101111111111;
    assign rom[3495]= 32'b00000000000010110100110111111111;
    assign rom[3496]= 32'b00000000000010110100111111111111;
    assign rom[3497]= 32'b00000000000010110101000111111111;
    assign rom[3498]= 32'b00000000000010110101001111111111;
    assign rom[3499]= 32'b00000000000010110101010111111111;
    assign rom[3500]= 32'b00000000000010110101011111111111;
    assign rom[3501]= 32'b00000000000010110101100111111111;
    assign rom[3502]= 32'b00000000000010110101101111111111;
    assign rom[3503]= 32'b00000000000010110101110111111111;
    assign rom[3504]= 32'b00000000000010110101111111111111;
    assign rom[3505]= 32'b00000000000010110110000111111111;
    assign rom[3506]= 32'b00000000000010110110001111111111;
    assign rom[3507]= 32'b00000000000010110110010111111111;
    assign rom[3508]= 32'b00000000000010110110011111111111;
    assign rom[3509]= 32'b00000000000010110110100111111111;
    assign rom[3510]= 32'b00000000000010110110101111111111;
    assign rom[3511]= 32'b00000000000010110110110111111111;
    assign rom[3512]= 32'b00000000000010110110111111111111;
    assign rom[3513]= 32'b00000000000010110111000111111111;
    assign rom[3514]= 32'b00000000000010110111001111111111;
    assign rom[3515]= 32'b00000000000010110111010111111111;
    assign rom[3516]= 32'b00000000000010110111011111111111;
    assign rom[3517]= 32'b00000000000010110111100111111111;
    assign rom[3518]= 32'b00000000000010110111101111111111;
    assign rom[3519]= 32'b00000000000010110111110111111111;
    assign rom[3520]= 32'b00000000000010110111111111111111;
    assign rom[3521]= 32'b00000000000010111000000111111111;
    assign rom[3522]= 32'b00000000000010111000001111111111;
    assign rom[3523]= 32'b00000000000010111000010111111111;
    assign rom[3524]= 32'b00000000000010111000011111111111;
    assign rom[3525]= 32'b00000000000010111000100111111111;
    assign rom[3526]= 32'b00000000000010111000101111111111;
    assign rom[3527]= 32'b00000000000010111000110111111111;
    assign rom[3528]= 32'b00000000000010111000111111111111;
    assign rom[3529]= 32'b00000000000010111001000111111111;
    assign rom[3530]= 32'b00000000000010111001001111111111;
    assign rom[3531]= 32'b00000000000010111001010111111111;
    assign rom[3532]= 32'b00000000000010111001011111111111;
    assign rom[3533]= 32'b00000000000010111001100111111111;
    assign rom[3534]= 32'b00000000000010111001101111111111;
    assign rom[3535]= 32'b00000000000010111001110111111111;
    assign rom[3536]= 32'b00000000000010111001111111111111;
    assign rom[3537]= 32'b00000000000010111010000111111111;
    assign rom[3538]= 32'b00000000000010111010001111111111;
    assign rom[3539]= 32'b00000000000010111010010111111111;
    assign rom[3540]= 32'b00000000000010111010011111111111;
    assign rom[3541]= 32'b00000000000010111010100111111111;
    assign rom[3542]= 32'b00000000000010111010101111111111;
    assign rom[3543]= 32'b00000000000010111010110111111111;
    assign rom[3544]= 32'b00000000000010111010111111111111;
    assign rom[3545]= 32'b00000000000010111011000111111111;
    assign rom[3546]= 32'b00000000000010111011001111111111;
    assign rom[3547]= 32'b00000000000010111011010111111111;
    assign rom[3548]= 32'b00000000000010111011011111111111;
    assign rom[3549]= 32'b00000000000010111011100111111111;
    assign rom[3550]= 32'b00000000000010111011101111111111;
    assign rom[3551]= 32'b00000000000010111011110111111111;
    assign rom[3552]= 32'b00000000000010111011111111111111;
    assign rom[3553]= 32'b00000000000010111100000111111111;
    assign rom[3554]= 32'b00000000000010111100001111111111;
    assign rom[3555]= 32'b00000000000010111100010111111111;
    assign rom[3556]= 32'b00000000000010111100011111111111;
    assign rom[3557]= 32'b00000000000010111100100111111111;
    assign rom[3558]= 32'b00000000000010111100101111111111;
    assign rom[3559]= 32'b00000000000010111100110111111111;
    assign rom[3560]= 32'b00000000000010111100111111111111;
    assign rom[3561]= 32'b00000000000010111101000111111111;
    assign rom[3562]= 32'b00000000000010111101001111111111;
    assign rom[3563]= 32'b00000000000010111101010111111111;
    assign rom[3564]= 32'b00000000000010111101011111111111;
    assign rom[3565]= 32'b00000000000010111101100111111111;
    assign rom[3566]= 32'b00000000000010111101101111111111;
    assign rom[3567]= 32'b00000000000010111101110111111111;
    assign rom[3568]= 32'b00000000000010111101111111111111;
    assign rom[3569]= 32'b00000000000010111110000111111111;
    assign rom[3570]= 32'b00000000000010111110001111111111;
    assign rom[3571]= 32'b00000000000010111110010111111111;
    assign rom[3572]= 32'b00000000000010111110011111111111;
    assign rom[3573]= 32'b00000000000010111110100111111111;
    assign rom[3574]= 32'b00000000000010111110101111111111;
    assign rom[3575]= 32'b00000000000010111110110111111111;
    assign rom[3576]= 32'b00000000000010111110111111111111;
    assign rom[3577]= 32'b00000000000010111111000111111111;
    assign rom[3578]= 32'b00000000000010111111001111111111;
    assign rom[3579]= 32'b00000000000010111111010111111111;
    assign rom[3580]= 32'b00000000000010111111011111111111;
    assign rom[3581]= 32'b00000000000010111111100111111111;
    assign rom[3582]= 32'b00000000000010111111101111111111;
    assign rom[3583]= 32'b00000000000010111111110111111111;
    assign rom[3584]= 32'b00000000000010111111111111111111;
    assign rom[3585]= 32'b00000000000011000000000111111111;
    assign rom[3586]= 32'b00000000000011000000001111111111;
    assign rom[3587]= 32'b00000000000011000000010111111111;
    assign rom[3588]= 32'b00000000000011000000011111111111;
    assign rom[3589]= 32'b00000000000011000000100111111111;
    assign rom[3590]= 32'b00000000000011000000101111111111;
    assign rom[3591]= 32'b00000000000011000000110111111111;
    assign rom[3592]= 32'b00000000000011000000111111111111;
    assign rom[3593]= 32'b00000000000011000001000111111111;
    assign rom[3594]= 32'b00000000000011000001001111111111;
    assign rom[3595]= 32'b00000000000011000001010111111111;
    assign rom[3596]= 32'b00000000000011000001011111111111;
    assign rom[3597]= 32'b00000000000011000001100111111111;
    assign rom[3598]= 32'b00000000000011000001101111111111;
    assign rom[3599]= 32'b00000000000011000001110111111111;
    assign rom[3600]= 32'b00000000000011000001111111111111;
    assign rom[3601]= 32'b00000000000011000010000111111111;
    assign rom[3602]= 32'b00000000000011000010001111111111;
    assign rom[3603]= 32'b00000000000011000010010111111111;
    assign rom[3604]= 32'b00000000000011000010011111111111;
    assign rom[3605]= 32'b00000000000011000010100111111111;
    assign rom[3606]= 32'b00000000000011000010101111111111;
    assign rom[3607]= 32'b00000000000011000010110111111111;
    assign rom[3608]= 32'b00000000000011000010111111111111;
    assign rom[3609]= 32'b00000000000011000011000111111111;
    assign rom[3610]= 32'b00000000000011000011001111111111;
    assign rom[3611]= 32'b00000000000011000011010111111111;
    assign rom[3612]= 32'b00000000000011000011011111111111;
    assign rom[3613]= 32'b00000000000011000011100111111111;
    assign rom[3614]= 32'b00000000000011000011101111111111;
    assign rom[3615]= 32'b00000000000011000011110111111111;
    assign rom[3616]= 32'b00000000000011000011111111111111;
    assign rom[3617]= 32'b00000000000011000100000111111111;
    assign rom[3618]= 32'b00000000000011000100001111111111;
    assign rom[3619]= 32'b00000000000011000100010111111111;
    assign rom[3620]= 32'b00000000000011000100011111111111;
    assign rom[3621]= 32'b00000000000011000100100111111111;
    assign rom[3622]= 32'b00000000000011000100101111111111;
    assign rom[3623]= 32'b00000000000011000100110111111111;
    assign rom[3624]= 32'b00000000000011000100111111111111;
    assign rom[3625]= 32'b00000000000011000101000111111111;
    assign rom[3626]= 32'b00000000000011000101001111111111;
    assign rom[3627]= 32'b00000000000011000101010111111111;
    assign rom[3628]= 32'b00000000000011000101011111111111;
    assign rom[3629]= 32'b00000000000011000101100111111111;
    assign rom[3630]= 32'b00000000000011000101101111111111;
    assign rom[3631]= 32'b00000000000011000101110111111111;
    assign rom[3632]= 32'b00000000000011000101111111111111;
    assign rom[3633]= 32'b00000000000011000110000111111111;
    assign rom[3634]= 32'b00000000000011000110001111111111;
    assign rom[3635]= 32'b00000000000011000110010111111111;
    assign rom[3636]= 32'b00000000000011000110011111111111;
    assign rom[3637]= 32'b00000000000011000110100111111111;
    assign rom[3638]= 32'b00000000000011000110101111111111;
    assign rom[3639]= 32'b00000000000011000110110111111111;
    assign rom[3640]= 32'b00000000000011000110111111111111;
    assign rom[3641]= 32'b00000000000011000111000111111111;
    assign rom[3642]= 32'b00000000000011000111001111111111;
    assign rom[3643]= 32'b00000000000011000111010111111111;
    assign rom[3644]= 32'b00000000000011000111011111111111;
    assign rom[3645]= 32'b00000000000011000111100111111111;
    assign rom[3646]= 32'b00000000000011000111101111111111;
    assign rom[3647]= 32'b00000000000011000111110111111111;
    assign rom[3648]= 32'b00000000000011000111111111111111;
    assign rom[3649]= 32'b00000000000011001000000111111111;
    assign rom[3650]= 32'b00000000000011001000001111111111;
    assign rom[3651]= 32'b00000000000011001000010111111111;
    assign rom[3652]= 32'b00000000000011001000011111111111;
    assign rom[3653]= 32'b00000000000011001000100111111111;
    assign rom[3654]= 32'b00000000000011001000101111111111;
    assign rom[3655]= 32'b00000000000011001000110111111111;
    assign rom[3656]= 32'b00000000000011001000111111111111;
    assign rom[3657]= 32'b00000000000011001001000111111111;
    assign rom[3658]= 32'b00000000000011001001001111111111;
    assign rom[3659]= 32'b00000000000011001001010111111111;
    assign rom[3660]= 32'b00000000000011001001011111111111;
    assign rom[3661]= 32'b00000000000011001001100111111111;
    assign rom[3662]= 32'b00000000000011001001101111111111;
    assign rom[3663]= 32'b00000000000011001001110111111111;
    assign rom[3664]= 32'b00000000000011001001111111111111;
    assign rom[3665]= 32'b00000000000011001010000111111111;
    assign rom[3666]= 32'b00000000000011001010001111111111;
    assign rom[3667]= 32'b00000000000011001010010111111111;
    assign rom[3668]= 32'b00000000000011001010011111111111;
    assign rom[3669]= 32'b00000000000011001010100111111111;
    assign rom[3670]= 32'b00000000000011001010101111111111;
    assign rom[3671]= 32'b00000000000011001010110111111111;
    assign rom[3672]= 32'b00000000000011001010111111111111;
    assign rom[3673]= 32'b00000000000011001011000111111111;
    assign rom[3674]= 32'b00000000000011001011001111111111;
    assign rom[3675]= 32'b00000000000011001011010111111111;
    assign rom[3676]= 32'b00000000000011001011011111111111;
    assign rom[3677]= 32'b00000000000011001011100111111111;
    assign rom[3678]= 32'b00000000000011001011101111111111;
    assign rom[3679]= 32'b00000000000011001011110111111111;
    assign rom[3680]= 32'b00000000000011001011111111111111;
    assign rom[3681]= 32'b00000000000011001100000111111111;
    assign rom[3682]= 32'b00000000000011001100001111111111;
    assign rom[3683]= 32'b00000000000011001100010111111111;
    assign rom[3684]= 32'b00000000000011001100011111111111;
    assign rom[3685]= 32'b00000000000011001100100111111111;
    assign rom[3686]= 32'b00000000000011001100101111111111;
    assign rom[3687]= 32'b00000000000011001100110111111111;
    assign rom[3688]= 32'b00000000000011001100111111111111;
    assign rom[3689]= 32'b00000000000011001101000111111111;
    assign rom[3690]= 32'b00000000000011001101001111111111;
    assign rom[3691]= 32'b00000000000011001101010111111111;
    assign rom[3692]= 32'b00000000000011001101011111111111;
    assign rom[3693]= 32'b00000000000011001101100111111111;
    assign rom[3694]= 32'b00000000000011001101101111111111;
    assign rom[3695]= 32'b00000000000011001101110111111111;
    assign rom[3696]= 32'b00000000000011001101111111111111;
    assign rom[3697]= 32'b00000000000011001110000111111111;
    assign rom[3698]= 32'b00000000000011001110001111111111;
    assign rom[3699]= 32'b00000000000011001110010111111111;
    assign rom[3700]= 32'b00000000000011001110011111111111;
    assign rom[3701]= 32'b00000000000011001110100111111111;
    assign rom[3702]= 32'b00000000000011001110101111111111;
    assign rom[3703]= 32'b00000000000011001110110111111111;
    assign rom[3704]= 32'b00000000000011001110111111111111;
    assign rom[3705]= 32'b00000000000011001111000111111111;
    assign rom[3706]= 32'b00000000000011001111001111111111;
    assign rom[3707]= 32'b00000000000011001111010111111111;
    assign rom[3708]= 32'b00000000000011001111011111111111;
    assign rom[3709]= 32'b00000000000011001111100111111111;
    assign rom[3710]= 32'b00000000000011001111101111111111;
    assign rom[3711]= 32'b00000000000011001111110111111111;
    assign rom[3712]= 32'b00000000000011001111111111111111;
    assign rom[3713]= 32'b00000000000011010000000111111111;
    assign rom[3714]= 32'b00000000000011010000001111111111;
    assign rom[3715]= 32'b00000000000011010000010111111111;
    assign rom[3716]= 32'b00000000000011010000011111111111;
    assign rom[3717]= 32'b00000000000011010000100111111111;
    assign rom[3718]= 32'b00000000000011010000101111111111;
    assign rom[3719]= 32'b00000000000011010000110111111111;
    assign rom[3720]= 32'b00000000000011010000111111111111;
    assign rom[3721]= 32'b00000000000011010001000111111111;
    assign rom[3722]= 32'b00000000000011010001001111111111;
    assign rom[3723]= 32'b00000000000011010001010111111111;
    assign rom[3724]= 32'b00000000000011010001011111111111;
    assign rom[3725]= 32'b00000000000011010001100111111111;
    assign rom[3726]= 32'b00000000000011010001101111111111;
    assign rom[3727]= 32'b00000000000011010001110111111111;
    assign rom[3728]= 32'b00000000000011010001111111111111;
    assign rom[3729]= 32'b00000000000011010010000111111111;
    assign rom[3730]= 32'b00000000000011010010001111111111;
    assign rom[3731]= 32'b00000000000011010010010111111111;
    assign rom[3732]= 32'b00000000000011010010011111111111;
    assign rom[3733]= 32'b00000000000011010010100111111111;
    assign rom[3734]= 32'b00000000000011010010101111111111;
    assign rom[3735]= 32'b00000000000011010010110111111111;
    assign rom[3736]= 32'b00000000000011010010111111111111;
    assign rom[3737]= 32'b00000000000011010011000111111111;
    assign rom[3738]= 32'b00000000000011010011001111111111;
    assign rom[3739]= 32'b00000000000011010011010111111111;
    assign rom[3740]= 32'b00000000000011010011011111111111;
    assign rom[3741]= 32'b00000000000011010011100111111111;
    assign rom[3742]= 32'b00000000000011010011101111111111;
    assign rom[3743]= 32'b00000000000011010011110111111111;
    assign rom[3744]= 32'b00000000000011010011111111111111;
    assign rom[3745]= 32'b00000000000011010100000111111111;
    assign rom[3746]= 32'b00000000000011010100001111111111;
    assign rom[3747]= 32'b00000000000011010100010111111111;
    assign rom[3748]= 32'b00000000000011010100011111111111;
    assign rom[3749]= 32'b00000000000011010100100111111111;
    assign rom[3750]= 32'b00000000000011010100101111111111;
    assign rom[3751]= 32'b00000000000011010100110111111111;
    assign rom[3752]= 32'b00000000000011010100111111111111;
    assign rom[3753]= 32'b00000000000011010101000111111111;
    assign rom[3754]= 32'b00000000000011010101001111111111;
    assign rom[3755]= 32'b00000000000011010101010111111111;
    assign rom[3756]= 32'b00000000000011010101011111111111;
    assign rom[3757]= 32'b00000000000011010101100111111111;
    assign rom[3758]= 32'b00000000000011010101101111111111;
    assign rom[3759]= 32'b00000000000011010101110111111111;
    assign rom[3760]= 32'b00000000000011010101111111111111;
    assign rom[3761]= 32'b00000000000011010110000111111111;
    assign rom[3762]= 32'b00000000000011010110001111111111;
    assign rom[3763]= 32'b00000000000011010110010111111111;
    assign rom[3764]= 32'b00000000000011010110011111111111;
    assign rom[3765]= 32'b00000000000011010110100111111111;
    assign rom[3766]= 32'b00000000000011010110101111111111;
    assign rom[3767]= 32'b00000000000011010110110111111111;
    assign rom[3768]= 32'b00000000000011010110111111111111;
    assign rom[3769]= 32'b00000000000011010111000111111111;
    assign rom[3770]= 32'b00000000000011010111001111111111;
    assign rom[3771]= 32'b00000000000011010111010111111111;
    assign rom[3772]= 32'b00000000000011010111011111111111;
    assign rom[3773]= 32'b00000000000011010111100111111111;
    assign rom[3774]= 32'b00000000000011010111101111111111;
    assign rom[3775]= 32'b00000000000011010111110111111111;
    assign rom[3776]= 32'b00000000000011010111111111111111;
    assign rom[3777]= 32'b00000000000011011000000111111111;
    assign rom[3778]= 32'b00000000000011011000001111111111;
    assign rom[3779]= 32'b00000000000011011000010111111111;
    assign rom[3780]= 32'b00000000000011011000011111111111;
    assign rom[3781]= 32'b00000000000011011000100111111111;
    assign rom[3782]= 32'b00000000000011011000101111111111;
    assign rom[3783]= 32'b00000000000011011000110111111111;
    assign rom[3784]= 32'b00000000000011011000111111111111;
    assign rom[3785]= 32'b00000000000011011001000111111111;
    assign rom[3786]= 32'b00000000000011011001001111111111;
    assign rom[3787]= 32'b00000000000011011001010111111111;
    assign rom[3788]= 32'b00000000000011011001011111111111;
    assign rom[3789]= 32'b00000000000011011001100111111111;
    assign rom[3790]= 32'b00000000000011011001101111111111;
    assign rom[3791]= 32'b00000000000011011001110111111111;
    assign rom[3792]= 32'b00000000000011011001111111111111;
    assign rom[3793]= 32'b00000000000011011010000111111111;
    assign rom[3794]= 32'b00000000000011011010001111111111;
    assign rom[3795]= 32'b00000000000011011010010111111111;
    assign rom[3796]= 32'b00000000000011011010011111111111;
    assign rom[3797]= 32'b00000000000011011010100111111111;
    assign rom[3798]= 32'b00000000000011011010101111111111;
    assign rom[3799]= 32'b00000000000011011010110111111111;
    assign rom[3800]= 32'b00000000000011011010111111111111;
    assign rom[3801]= 32'b00000000000011011011000111111111;
    assign rom[3802]= 32'b00000000000011011011001111111111;
    assign rom[3803]= 32'b00000000000011011011010111111111;
    assign rom[3804]= 32'b00000000000011011011011111111111;
    assign rom[3805]= 32'b00000000000011011011100111111111;
    assign rom[3806]= 32'b00000000000011011011101111111111;
    assign rom[3807]= 32'b00000000000011011011110111111111;
    assign rom[3808]= 32'b00000000000011011011111111111111;
    assign rom[3809]= 32'b00000000000011011100000111111111;
    assign rom[3810]= 32'b00000000000011011100001111111111;
    assign rom[3811]= 32'b00000000000011011100010111111111;
    assign rom[3812]= 32'b00000000000011011100011111111111;
    assign rom[3813]= 32'b00000000000011011100100111111111;
    assign rom[3814]= 32'b00000000000011011100101111111111;
    assign rom[3815]= 32'b00000000000011011100110111111111;
    assign rom[3816]= 32'b00000000000011011100111111111111;
    assign rom[3817]= 32'b00000000000011011101000111111111;
    assign rom[3818]= 32'b00000000000011011101001111111111;
    assign rom[3819]= 32'b00000000000011011101010111111111;
    assign rom[3820]= 32'b00000000000011011101011111111111;
    assign rom[3821]= 32'b00000000000011011101100111111111;
    assign rom[3822]= 32'b00000000000011011101101111111111;
    assign rom[3823]= 32'b00000000000011011101110111111111;
    assign rom[3824]= 32'b00000000000011011101111111111111;
    assign rom[3825]= 32'b00000000000011011110000111111111;
    assign rom[3826]= 32'b00000000000011011110001111111111;
    assign rom[3827]= 32'b00000000000011011110010111111111;
    assign rom[3828]= 32'b00000000000011011110011111111111;
    assign rom[3829]= 32'b00000000000011011110100111111111;
    assign rom[3830]= 32'b00000000000011011110101111111111;
    assign rom[3831]= 32'b00000000000011011110110111111111;
    assign rom[3832]= 32'b00000000000011011110111111111111;
    assign rom[3833]= 32'b00000000000011011111000111111111;
    assign rom[3834]= 32'b00000000000011011111001111111111;
    assign rom[3835]= 32'b00000000000011011111010111111111;
    assign rom[3836]= 32'b00000000000011011111011111111111;
    assign rom[3837]= 32'b00000000000011011111100111111111;
    assign rom[3838]= 32'b00000000000011011111101111111111;
    assign rom[3839]= 32'b00000000000011011111110111111111;
    assign rom[3840]= 32'b00000000000011011111111111111111;
    assign rom[3841]= 32'b00000000000011100000000111111111;
    assign rom[3842]= 32'b00000000000011100000001111111111;
    assign rom[3843]= 32'b00000000000011100000010111111111;
    assign rom[3844]= 32'b00000000000011100000011111111111;
    assign rom[3845]= 32'b00000000000011100000100111111111;
    assign rom[3846]= 32'b00000000000011100000101111111111;
    assign rom[3847]= 32'b00000000000011100000110111111111;
    assign rom[3848]= 32'b00000000000011100000111111111111;
    assign rom[3849]= 32'b00000000000011100001000111111111;
    assign rom[3850]= 32'b00000000000011100001001111111111;
    assign rom[3851]= 32'b00000000000011100001010111111111;
    assign rom[3852]= 32'b00000000000011100001011111111111;
    assign rom[3853]= 32'b00000000000011100001100111111111;
    assign rom[3854]= 32'b00000000000011100001101111111111;
    assign rom[3855]= 32'b00000000000011100001110111111111;
    assign rom[3856]= 32'b00000000000011100001111111111111;
    assign rom[3857]= 32'b00000000000011100010000111111111;
    assign rom[3858]= 32'b00000000000011100010001111111111;
    assign rom[3859]= 32'b00000000000011100010010111111111;
    assign rom[3860]= 32'b00000000000011100010011111111111;
    assign rom[3861]= 32'b00000000000011100010100111111111;
    assign rom[3862]= 32'b00000000000011100010101111111111;
    assign rom[3863]= 32'b00000000000011100010110111111111;
    assign rom[3864]= 32'b00000000000011100010111111111111;
    assign rom[3865]= 32'b00000000000011100011000111111111;
    assign rom[3866]= 32'b00000000000011100011001111111111;
    assign rom[3867]= 32'b00000000000011100011010111111111;
    assign rom[3868]= 32'b00000000000011100011011111111111;
    assign rom[3869]= 32'b00000000000011100011100111111111;
    assign rom[3870]= 32'b00000000000011100011101111111111;
    assign rom[3871]= 32'b00000000000011100011110111111111;
    assign rom[3872]= 32'b00000000000011100011111111111111;
    assign rom[3873]= 32'b00000000000011100100000111111111;
    assign rom[3874]= 32'b00000000000011100100001111111111;
    assign rom[3875]= 32'b00000000000011100100010111111111;
    assign rom[3876]= 32'b00000000000011100100011111111111;
    assign rom[3877]= 32'b00000000000011100100100111111111;
    assign rom[3878]= 32'b00000000000011100100101111111111;
    assign rom[3879]= 32'b00000000000011100100110111111111;
    assign rom[3880]= 32'b00000000000011100100111111111111;
    assign rom[3881]= 32'b00000000000011100101000111111111;
    assign rom[3882]= 32'b00000000000011100101001111111111;
    assign rom[3883]= 32'b00000000000011100101010111111111;
    assign rom[3884]= 32'b00000000000011100101011111111111;
    assign rom[3885]= 32'b00000000000011100101100111111111;
    assign rom[3886]= 32'b00000000000011100101101111111111;
    assign rom[3887]= 32'b00000000000011100101110111111111;
    assign rom[3888]= 32'b00000000000011100101111111111111;
    assign rom[3889]= 32'b00000000000011100110000111111111;
    assign rom[3890]= 32'b00000000000011100110001111111111;
    assign rom[3891]= 32'b00000000000011100110010111111111;
    assign rom[3892]= 32'b00000000000011100110011111111111;
    assign rom[3893]= 32'b00000000000011100110100111111111;
    assign rom[3894]= 32'b00000000000011100110101111111111;
    assign rom[3895]= 32'b00000000000011100110110111111111;
    assign rom[3896]= 32'b00000000000011100110111111111111;
    assign rom[3897]= 32'b00000000000011100111000111111111;
    assign rom[3898]= 32'b00000000000011100111001111111111;
    assign rom[3899]= 32'b00000000000011100111010111111111;
    assign rom[3900]= 32'b00000000000011100111011111111111;
    assign rom[3901]= 32'b00000000000011100111100111111111;
    assign rom[3902]= 32'b00000000000011100111101111111111;
    assign rom[3903]= 32'b00000000000011100111110111111111;
    assign rom[3904]= 32'b00000000000011100111111111111111;
    assign rom[3905]= 32'b00000000000011101000000111111111;
    assign rom[3906]= 32'b00000000000011101000001111111111;
    assign rom[3907]= 32'b00000000000011101000010111111111;
    assign rom[3908]= 32'b00000000000011101000011111111111;
    assign rom[3909]= 32'b00000000000011101000100111111111;
    assign rom[3910]= 32'b00000000000011101000101111111111;
    assign rom[3911]= 32'b00000000000011101000110111111111;
    assign rom[3912]= 32'b00000000000011101000111111111111;
    assign rom[3913]= 32'b00000000000011101001000111111111;
    assign rom[3914]= 32'b00000000000011101001001111111111;
    assign rom[3915]= 32'b00000000000011101001010111111111;
    assign rom[3916]= 32'b00000000000011101001011111111111;
    assign rom[3917]= 32'b00000000000011101001100111111111;
    assign rom[3918]= 32'b00000000000011101001101111111111;
    assign rom[3919]= 32'b00000000000011101001110111111111;
    assign rom[3920]= 32'b00000000000011101001111111111111;
    assign rom[3921]= 32'b00000000000011101010000111111111;
    assign rom[3922]= 32'b00000000000011101010001111111111;
    assign rom[3923]= 32'b00000000000011101010010111111111;
    assign rom[3924]= 32'b00000000000011101010011111111111;
    assign rom[3925]= 32'b00000000000011101010100111111111;
    assign rom[3926]= 32'b00000000000011101010101111111111;
    assign rom[3927]= 32'b00000000000011101010110111111111;
    assign rom[3928]= 32'b00000000000011101010111111111111;
    assign rom[3929]= 32'b00000000000011101011000111111111;
    assign rom[3930]= 32'b00000000000011101011001111111111;
    assign rom[3931]= 32'b00000000000011101011010111111111;
    assign rom[3932]= 32'b00000000000011101011011111111111;
    assign rom[3933]= 32'b00000000000011101011100111111111;
    assign rom[3934]= 32'b00000000000011101011101111111111;
    assign rom[3935]= 32'b00000000000011101011110111111111;
    assign rom[3936]= 32'b00000000000011101011111111111111;
    assign rom[3937]= 32'b00000000000011101100000111111111;
    assign rom[3938]= 32'b00000000000011101100001111111111;
    assign rom[3939]= 32'b00000000000011101100010111111111;
    assign rom[3940]= 32'b00000000000011101100011111111111;
    assign rom[3941]= 32'b00000000000011101100100111111111;
    assign rom[3942]= 32'b00000000000011101100101111111111;
    assign rom[3943]= 32'b00000000000011101100110111111111;
    assign rom[3944]= 32'b00000000000011101100111111111111;
    assign rom[3945]= 32'b00000000000011101101000111111111;
    assign rom[3946]= 32'b00000000000011101101001111111111;
    assign rom[3947]= 32'b00000000000011101101010111111111;
    assign rom[3948]= 32'b00000000000011101101011111111111;
    assign rom[3949]= 32'b00000000000011101101100111111111;
    assign rom[3950]= 32'b00000000000011101101101111111111;
    assign rom[3951]= 32'b00000000000011101101110111111111;
    assign rom[3952]= 32'b00000000000011101101111111111111;
    assign rom[3953]= 32'b00000000000011101110000111111111;
    assign rom[3954]= 32'b00000000000011101110001111111111;
    assign rom[3955]= 32'b00000000000011101110010111111111;
    assign rom[3956]= 32'b00000000000011101110011111111111;
    assign rom[3957]= 32'b00000000000011101110100111111111;
    assign rom[3958]= 32'b00000000000011101110101111111111;
    assign rom[3959]= 32'b00000000000011101110110111111111;
    assign rom[3960]= 32'b00000000000011101110111111111111;
    assign rom[3961]= 32'b00000000000011101111000111111111;
    assign rom[3962]= 32'b00000000000011101111001111111111;
    assign rom[3963]= 32'b00000000000011101111010111111111;
    assign rom[3964]= 32'b00000000000011101111011111111111;
    assign rom[3965]= 32'b00000000000011101111100111111111;
    assign rom[3966]= 32'b00000000000011101111101111111111;
    assign rom[3967]= 32'b00000000000011101111110111111111;
    assign rom[3968]= 32'b00000000000011101111111111111111;
    assign rom[3969]= 32'b00000000000011110000000111111111;
    assign rom[3970]= 32'b00000000000011110000001111111111;
    assign rom[3971]= 32'b00000000000011110000010111111111;
    assign rom[3972]= 32'b00000000000011110000011111111111;
    assign rom[3973]= 32'b00000000000011110000100111111111;
    assign rom[3974]= 32'b00000000000011110000101111111111;
    assign rom[3975]= 32'b00000000000011110000110111111111;
    assign rom[3976]= 32'b00000000000011110000111111111111;
    assign rom[3977]= 32'b00000000000011110001000111111111;
    assign rom[3978]= 32'b00000000000011110001001111111111;
    assign rom[3979]= 32'b00000000000011110001010111111111;
    assign rom[3980]= 32'b00000000000011110001011111111111;
    assign rom[3981]= 32'b00000000000011110001100111111111;
    assign rom[3982]= 32'b00000000000011110001101111111111;
    assign rom[3983]= 32'b00000000000011110001110111111111;
    assign rom[3984]= 32'b00000000000011110001111111111111;
    assign rom[3985]= 32'b00000000000011110010000111111111;
    assign rom[3986]= 32'b00000000000011110010001111111111;
    assign rom[3987]= 32'b00000000000011110010010111111111;
    assign rom[3988]= 32'b00000000000011110010011111111111;
    assign rom[3989]= 32'b00000000000011110010100111111111;
    assign rom[3990]= 32'b00000000000011110010101111111111;
    assign rom[3991]= 32'b00000000000011110010110111111111;
    assign rom[3992]= 32'b00000000000011110010111111111111;
    assign rom[3993]= 32'b00000000000011110011000111111111;
    assign rom[3994]= 32'b00000000000011110011001111111111;
    assign rom[3995]= 32'b00000000000011110011010111111111;
    assign rom[3996]= 32'b00000000000011110011011111111111;
    assign rom[3997]= 32'b00000000000011110011100111111111;
    assign rom[3998]= 32'b00000000000011110011101111111111;
    assign rom[3999]= 32'b00000000000011110011110111111111;
    assign rom[4000]= 32'b00000000000011110011111111111111;
    assign rom[4001]= 32'b00000000000011110100000111111111;
    assign rom[4002]= 32'b00000000000011110100001111111111;
    assign rom[4003]= 32'b00000000000011110100010111111111;
    assign rom[4004]= 32'b00000000000011110100011111111111;
    assign rom[4005]= 32'b00000000000011110100100111111111;
    assign rom[4006]= 32'b00000000000011110100101111111111;
    assign rom[4007]= 32'b00000000000011110100110111111111;
    assign rom[4008]= 32'b00000000000011110100111111111111;
    assign rom[4009]= 32'b00000000000011110101000111111111;
    assign rom[4010]= 32'b00000000000011110101001111111111;
    assign rom[4011]= 32'b00000000000011110101010111111111;
    assign rom[4012]= 32'b00000000000011110101011111111111;
    assign rom[4013]= 32'b00000000000011110101100111111111;
    assign rom[4014]= 32'b00000000000011110101101111111111;
    assign rom[4015]= 32'b00000000000011110101110111111111;
    assign rom[4016]= 32'b00000000000011110101111111111111;
    assign rom[4017]= 32'b00000000000011110110000111111111;
    assign rom[4018]= 32'b00000000000011110110001111111111;
    assign rom[4019]= 32'b00000000000011110110010111111111;
    assign rom[4020]= 32'b00000000000011110110011111111111;
    assign rom[4021]= 32'b00000000000011110110100111111111;
    assign rom[4022]= 32'b00000000000011110110101111111111;
    assign rom[4023]= 32'b00000000000011110110110111111111;
    assign rom[4024]= 32'b00000000000011110110111111111111;
    assign rom[4025]= 32'b00000000000011110111000111111111;
    assign rom[4026]= 32'b00000000000011110111001111111111;
    assign rom[4027]= 32'b00000000000011110111010111111111;
    assign rom[4028]= 32'b00000000000011110111011111111111;
    assign rom[4029]= 32'b00000000000011110111100111111111;
    assign rom[4030]= 32'b00000000000011110111101111111111;
    assign rom[4031]= 32'b00000000000011110111110111111111;
    assign rom[4032]= 32'b00000000000011110111111111111111;
    assign rom[4033]= 32'b00000000000011111000000111111111;
    assign rom[4034]= 32'b00000000000011111000001111111111;
    assign rom[4035]= 32'b00000000000011111000010111111111;
    assign rom[4036]= 32'b00000000000011111000011111111111;
    assign rom[4037]= 32'b00000000000011111000100111111111;
    assign rom[4038]= 32'b00000000000011111000101111111111;
    assign rom[4039]= 32'b00000000000011111000110111111111;
    assign rom[4040]= 32'b00000000000011111000111111111111;
    assign rom[4041]= 32'b00000000000011111001000111111111;
    assign rom[4042]= 32'b00000000000011111001001111111111;
    assign rom[4043]= 32'b00000000000011111001010111111111;
    assign rom[4044]= 32'b00000000000011111001011111111111;
    assign rom[4045]= 32'b00000000000011111001100111111111;
    assign rom[4046]= 32'b00000000000011111001101111111111;
    assign rom[4047]= 32'b00000000000011111001110111111111;
    assign rom[4048]= 32'b00000000000011111001111111111111;
    assign rom[4049]= 32'b00000000000011111010000111111111;
    assign rom[4050]= 32'b00000000000011111010001111111111;
    assign rom[4051]= 32'b00000000000011111010010111111111;
    assign rom[4052]= 32'b00000000000011111010011111111111;
    assign rom[4053]= 32'b00000000000011111010100111111111;
    assign rom[4054]= 32'b00000000000011111010101111111111;
    assign rom[4055]= 32'b00000000000011111010110111111111;
    assign rom[4056]= 32'b00000000000011111010111111111111;
    assign rom[4057]= 32'b00000000000011111011000111111111;
    assign rom[4058]= 32'b00000000000011111011001111111111;
    assign rom[4059]= 32'b00000000000011111011010111111111;
    assign rom[4060]= 32'b00000000000011111011011111111111;
    assign rom[4061]= 32'b00000000000011111011100111111111;
    assign rom[4062]= 32'b00000000000011111011101111111111;
    assign rom[4063]= 32'b00000000000011111011110111111111;
    assign rom[4064]= 32'b00000000000011111011111111111111;
    assign rom[4065]= 32'b00000000000011111100000111111111;
    assign rom[4066]= 32'b00000000000011111100001111111111;
    assign rom[4067]= 32'b00000000000011111100010111111111;
    assign rom[4068]= 32'b00000000000011111100011111111111;
    assign rom[4069]= 32'b00000000000011111100100111111111;
    assign rom[4070]= 32'b00000000000011111100101111111111;
    assign rom[4071]= 32'b00000000000011111100110111111111;
    assign rom[4072]= 32'b00000000000011111100111111111111;
    assign rom[4073]= 32'b00000000000011111101000111111111;
    assign rom[4074]= 32'b00000000000011111101001111111111;
    assign rom[4075]= 32'b00000000000011111101010111111111;
    assign rom[4076]= 32'b00000000000011111101011111111111;
    assign rom[4077]= 32'b00000000000011111101100111111111;
    assign rom[4078]= 32'b00000000000011111101101111111111;
    assign rom[4079]= 32'b00000000000011111101110111111111;
    assign rom[4080]= 32'b00000000000011111101111111111111;
    assign rom[4081]= 32'b00000000000011111110000111111111;
    assign rom[4082]= 32'b00000000000011111110001111111111;
    assign rom[4083]= 32'b00000000000011111110010111111111;
    assign rom[4084]= 32'b00000000000011111110011111111111;
    assign rom[4085]= 32'b00000000000011111110100111111111;
    assign rom[4086]= 32'b00000000000011111110101111111111;
    assign rom[4087]= 32'b00000000000011111110110111111111;
    assign rom[4088]= 32'b00000000000011111110111111111111;
    assign rom[4089]= 32'b00000000000011111111000111111111;
    assign rom[4090]= 32'b00000000000011111111001111111111;
    assign rom[4091]= 32'b00000000000011111111010111111111;
    assign rom[4092]= 32'b00000000000011111111011111111111;
    assign rom[4093]= 32'b00000000000011111111100111111111;
    assign rom[4094]= 32'b00000000000011111111101111111111;
    assign rom[4095]= 32'b00000000000011111111110111111111;


    always @(*) begin
        data_out = rom[addr];
    end
endmodule
